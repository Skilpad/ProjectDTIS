
module reg_0 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n142, n350, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n538, n539, n540, n542,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  DF3 Dout_reg_31_ ( .D(n560), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n561), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n562), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n563), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n564), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n565), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n566), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n567), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n568), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n569), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n570), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n571), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n572), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n573), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n574), .C(Clk), .Q(Dout[17]), .QN(n548) );
  DF3 Dout_reg_16_ ( .D(n575), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_15_ ( .D(n576), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n577), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_13_ ( .D(n578), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_12_ ( .D(n579), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_11_ ( .D(n580), .C(Clk), .Q(n142) );
  DF3 Dout_reg_10_ ( .D(n581), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_9_ ( .D(n582), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_8_ ( .D(n583), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_7_ ( .D(n584), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_6_ ( .D(n585), .C(Clk), .Q(Dout[6]), .QN(n544) );
  DF3 Dout_reg_5_ ( .D(n586), .C(Clk), .Q(Dout[5]), .QN(n538) );
  DF3 Dout_reg_4_ ( .D(n587), .C(Clk), .Q(Dout[4]), .QN(n546) );
  DF3 Dout_reg_3_ ( .D(n588), .C(Clk), .Q(n350) );
  DF3 Dout_reg_2_ ( .D(n589), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_1_ ( .D(n590), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_0_ ( .D(n591), .C(Clk), .Q(Dout[0]) );
  INV3 U3 ( .A(n538), .Q(n539) );
  CLKIN6 U4 ( .A(n142), .Q(n540) );
  INV12 U5 ( .A(n540), .Q(Dout[11]) );
  INV3 U6 ( .A(n350), .Q(n542) );
  INV6 U7 ( .A(n542), .Q(Dout[3]) );
  INV3 U8 ( .A(n544), .Q(n545) );
  INV3 U9 ( .A(n546), .Q(n547) );
  INV3 U10 ( .A(n548), .Q(n549) );
  AOI220 U11 ( .A(Din[28]), .B(n559), .C(n553), .D(Dout[28]), .Q(n38) );
  INV3 U12 ( .A(n558), .Q(n559) );
  CLKBU2 U13 ( .A(n550), .Q(n552) );
  CLKBU2 U14 ( .A(n550), .Q(n553) );
  CLKBU2 U15 ( .A(n35), .Q(n556) );
  CLKBU2 U16 ( .A(n35), .Q(n557) );
  CLKBU2 U17 ( .A(n551), .Q(n554) );
  CLKBU2 U18 ( .A(n551), .Q(n555) );
  INV3 U19 ( .A(n62), .Q(n587) );
  INV3 U20 ( .A(n61), .Q(n586) );
  INV3 U21 ( .A(n60), .Q(n585) );
  INV3 U22 ( .A(n59), .Q(n584) );
  INV3 U23 ( .A(n58), .Q(n583) );
  INV3 U24 ( .A(n57), .Q(n582) );
  INV3 U25 ( .A(n56), .Q(n581) );
  INV3 U26 ( .A(n53), .Q(n578) );
  INV3 U27 ( .A(n52), .Q(n577) );
  INV3 U28 ( .A(n50), .Q(n575) );
  INV3 U29 ( .A(n49), .Q(n574) );
  INV3 U30 ( .A(n48), .Q(n573) );
  INV3 U31 ( .A(n47), .Q(n572) );
  INV3 U32 ( .A(n45), .Q(n570) );
  NOR20 U33 ( .A(Load), .B(Reset), .Q(n550) );
  NOR20 U34 ( .A(Load), .B(Reset), .Q(n551) );
  NOR20 U35 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U36 ( .A(n34), .Q(n558) );
  NOR21 U37 ( .A(n552), .B(Reset), .Q(n34) );
  INV3 U38 ( .A(n66), .Q(n591) );
  AOI220 U39 ( .A(Din[0]), .B(n559), .C(n552), .D(Dout[0]), .Q(n66) );
  INV3 U40 ( .A(n65), .Q(n590) );
  AOI220 U41 ( .A(Din[1]), .B(n34), .C(n553), .D(Dout[1]), .Q(n65) );
  INV3 U42 ( .A(n64), .Q(n589) );
  AOI220 U43 ( .A(Din[2]), .B(n559), .C(n553), .D(Dout[2]), .Q(n64) );
  INV3 U44 ( .A(n63), .Q(n588) );
  AOI220 U45 ( .A(Din[3]), .B(n34), .C(n552), .D(Dout[3]), .Q(n63) );
  INV3 U46 ( .A(n55), .Q(n580) );
  AOI220 U47 ( .A(Din[11]), .B(n34), .C(n557), .D(Dout[11]), .Q(n55) );
  INV3 U48 ( .A(n54), .Q(n579) );
  AOI220 U49 ( .A(Din[12]), .B(n559), .C(n556), .D(Dout[12]), .Q(n54) );
  INV3 U50 ( .A(n51), .Q(n576) );
  AOI220 U51 ( .A(Din[15]), .B(n34), .C(n552), .D(Dout[15]), .Q(n51) );
  INV3 U52 ( .A(n46), .Q(n571) );
  AOI220 U53 ( .A(Din[20]), .B(n559), .C(n556), .D(Dout[20]), .Q(n46) );
  INV3 U54 ( .A(n44), .Q(n569) );
  AOI220 U55 ( .A(Din[22]), .B(n559), .C(n556), .D(Dout[22]), .Q(n44) );
  INV3 U56 ( .A(n43), .Q(n568) );
  AOI220 U57 ( .A(Din[23]), .B(n34), .C(n557), .D(Dout[23]), .Q(n43) );
  INV3 U58 ( .A(n42), .Q(n567) );
  AOI220 U59 ( .A(Din[24]), .B(n559), .C(n554), .D(Dout[24]), .Q(n42) );
  INV3 U60 ( .A(n41), .Q(n566) );
  AOI220 U61 ( .A(Din[25]), .B(n34), .C(n555), .D(Dout[25]), .Q(n41) );
  INV3 U62 ( .A(n40), .Q(n565) );
  AOI220 U63 ( .A(Din[26]), .B(n559), .C(n557), .D(Dout[26]), .Q(n40) );
  INV3 U64 ( .A(n39), .Q(n564) );
  AOI220 U65 ( .A(Din[27]), .B(n34), .C(n552), .D(Dout[27]), .Q(n39) );
  INV3 U66 ( .A(n38), .Q(n563) );
  INV3 U67 ( .A(n37), .Q(n562) );
  AOI220 U68 ( .A(Din[29]), .B(n34), .C(n554), .D(Dout[29]), .Q(n37) );
  INV3 U69 ( .A(n36), .Q(n561) );
  AOI221 U70 ( .A(Din[30]), .B(n559), .C(n556), .D(Dout[30]), .Q(n36) );
  INV3 U71 ( .A(n33), .Q(n560) );
  AOI221 U72 ( .A(Din[31]), .B(n34), .C(n557), .D(Dout[31]), .Q(n33) );
  AOI220 U73 ( .A(Din[14]), .B(n559), .C(n555), .D(Dout[14]), .Q(n52) );
  AOI220 U74 ( .A(Din[9]), .B(n34), .C(n555), .D(Dout[9]), .Q(n57) );
  AOI220 U75 ( .A(Din[16]), .B(n559), .C(n553), .D(Dout[16]), .Q(n50) );
  AOI220 U76 ( .A(Din[21]), .B(n34), .C(n555), .D(Dout[21]), .Q(n45) );
  AOI220 U77 ( .A(Din[7]), .B(n34), .C(n555), .D(Dout[7]), .Q(n59) );
  AOI220 U78 ( .A(Din[4]), .B(n559), .C(n553), .D(n547), .Q(n62) );
  AOI220 U79 ( .A(Din[19]), .B(n34), .C(n553), .D(Dout[19]), .Q(n47) );
  AOI220 U80 ( .A(Din[13]), .B(n34), .C(n557), .D(Dout[13]), .Q(n53) );
  AOI220 U81 ( .A(Din[8]), .B(n559), .C(n554), .D(Dout[8]), .Q(n58) );
  AOI220 U82 ( .A(Din[10]), .B(n559), .C(n556), .D(Dout[10]), .Q(n56) );
  AOI220 U83 ( .A(Din[6]), .B(n559), .C(n554), .D(n545), .Q(n60) );
  AOI220 U84 ( .A(Din[18]), .B(n559), .C(n552), .D(Dout[18]), .Q(n48) );
  AOI220 U85 ( .A(Din[5]), .B(n34), .C(n539), .D(n554), .Q(n61) );
  AOI220 U86 ( .A(Din[17]), .B(n559), .C(n554), .D(n549), .Q(n49) );
endmodule


module reg_33 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504;

  DF3 Dout_reg_31_ ( .D(n473), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n474), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n475), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n476), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n477), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n478), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n479), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n480), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n481), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n482), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n483), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n484), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n485), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n486), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n487), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_16_ ( .D(n488), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_13_ ( .D(n489), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_12_ ( .D(n490), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_6_ ( .D(n491), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_9_ ( .D(n492), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_7_ ( .D(n493), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_1_ ( .D(n494), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_4_ ( .D(n496), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_0_ ( .D(n497), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_10_ ( .D(n498), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_15_ ( .D(n499), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n500), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_8_ ( .D(n502), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_3_ ( .D(n503), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_2_ ( .D(n504), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_11_ ( .D(n495), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_5_ ( .D(n501), .C(Clk), .Q(Dout[5]) );
  AOI220 U3 ( .A(Din[28]), .B(n472), .C(n466), .D(Dout[28]), .Q(n38) );
  INV3 U4 ( .A(n471), .Q(n472) );
  CLKBU2 U5 ( .A(n463), .Q(n465) );
  CLKBU2 U6 ( .A(n464), .Q(n467) );
  CLKBU2 U7 ( .A(n464), .Q(n468) );
  CLKBU2 U8 ( .A(n35), .Q(n469) );
  CLKBU2 U9 ( .A(n35), .Q(n470) );
  CLKBU2 U10 ( .A(n463), .Q(n466) );
  INV3 U11 ( .A(n63), .Q(n501) );
  INV3 U12 ( .A(n66), .Q(n504) );
  INV3 U13 ( .A(n65), .Q(n503) );
  INV3 U14 ( .A(n64), .Q(n502) );
  INV3 U15 ( .A(n62), .Q(n500) );
  INV3 U16 ( .A(n60), .Q(n498) );
  INV3 U17 ( .A(n58), .Q(n496) );
  INV3 U18 ( .A(n56), .Q(n494) );
  INV3 U19 ( .A(n55), .Q(n493) );
  INV3 U20 ( .A(n54), .Q(n492) );
  INV3 U21 ( .A(n53), .Q(n491) );
  INV3 U22 ( .A(n51), .Q(n489) );
  INV3 U23 ( .A(n50), .Q(n488) );
  INV3 U24 ( .A(n49), .Q(n487) );
  INV3 U25 ( .A(n48), .Q(n486) );
  INV3 U26 ( .A(n47), .Q(n485) );
  INV3 U27 ( .A(n45), .Q(n483) );
  INV3 U28 ( .A(n59), .Q(n497) );
  AOI220 U29 ( .A(Din[0]), .B(n34), .C(n468), .D(Dout[0]), .Q(n59) );
  INV3 U30 ( .A(n43), .Q(n481) );
  AOI220 U31 ( .A(Din[23]), .B(n34), .C(n470), .D(Dout[23]), .Q(n43) );
  INV3 U32 ( .A(n40), .Q(n478) );
  AOI220 U33 ( .A(Din[26]), .B(n472), .C(n470), .D(Dout[26]), .Q(n40) );
  INV3 U34 ( .A(n44), .Q(n482) );
  AOI220 U35 ( .A(Din[22]), .B(n472), .C(n469), .D(Dout[22]), .Q(n44) );
  INV3 U36 ( .A(n42), .Q(n480) );
  AOI220 U37 ( .A(Din[24]), .B(n472), .C(n467), .D(Dout[24]), .Q(n42) );
  INV3 U38 ( .A(n57), .Q(n495) );
  AOI220 U39 ( .A(Din[11]), .B(n34), .C(n468), .D(Dout[11]), .Q(n57) );
  INV3 U40 ( .A(n41), .Q(n479) );
  AOI220 U41 ( .A(Din[25]), .B(n34), .C(n468), .D(Dout[25]), .Q(n41) );
  INV3 U42 ( .A(n39), .Q(n477) );
  AOI220 U43 ( .A(Din[27]), .B(n34), .C(n465), .D(Dout[27]), .Q(n39) );
  INV3 U44 ( .A(n52), .Q(n490) );
  AOI220 U45 ( .A(Din[12]), .B(n472), .C(n468), .D(Dout[12]), .Q(n52) );
  INV3 U46 ( .A(n38), .Q(n476) );
  INV3 U47 ( .A(n37), .Q(n475) );
  AOI220 U48 ( .A(Din[29]), .B(n34), .C(n467), .D(Dout[29]), .Q(n37) );
  INV3 U49 ( .A(n33), .Q(n473) );
  AOI221 U50 ( .A(Din[31]), .B(n34), .C(n470), .D(Dout[31]), .Q(n33) );
  INV3 U51 ( .A(n46), .Q(n484) );
  AOI220 U52 ( .A(Din[20]), .B(n472), .C(n469), .D(Dout[20]), .Q(n46) );
  INV3 U53 ( .A(n36), .Q(n474) );
  AOI221 U54 ( .A(Din[30]), .B(n472), .C(n469), .D(Dout[30]), .Q(n36) );
  INV3 U55 ( .A(n61), .Q(n499) );
  AOI220 U56 ( .A(Din[15]), .B(n34), .C(n467), .D(Dout[15]), .Q(n61) );
  NOR20 U57 ( .A(Load), .B(Reset), .Q(n463) );
  NOR20 U58 ( .A(Load), .B(Reset), .Q(n464) );
  NOR20 U59 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U60 ( .A(n34), .Q(n471) );
  NOR21 U61 ( .A(n465), .B(Reset), .Q(n34) );
  AOI220 U62 ( .A(Din[1]), .B(n472), .C(n469), .D(Dout[1]), .Q(n56) );
  AOI220 U63 ( .A(Din[14]), .B(n472), .C(n466), .D(Dout[14]), .Q(n62) );
  AOI220 U64 ( .A(Din[9]), .B(n472), .C(n469), .D(Dout[9]), .Q(n54) );
  AOI220 U65 ( .A(Din[16]), .B(n472), .C(n466), .D(Dout[16]), .Q(n50) );
  AOI220 U66 ( .A(Din[21]), .B(n34), .C(n468), .D(Dout[21]), .Q(n45) );
  AOI220 U67 ( .A(Din[7]), .B(n34), .C(n470), .D(Dout[7]), .Q(n55) );
  AOI220 U68 ( .A(Din[4]), .B(n472), .C(n467), .D(Dout[4]), .Q(n58) );
  AOI220 U69 ( .A(Din[19]), .B(n34), .C(n466), .D(Dout[19]), .Q(n47) );
  AOI220 U70 ( .A(Din[2]), .B(n472), .C(n465), .D(Dout[2]), .Q(n66) );
  AOI220 U71 ( .A(Din[13]), .B(n34), .C(n465), .D(Dout[13]), .Q(n51) );
  AOI220 U72 ( .A(Din[8]), .B(n472), .C(n466), .D(Dout[8]), .Q(n64) );
  AOI220 U73 ( .A(Din[10]), .B(n472), .C(n467), .D(Dout[10]), .Q(n60) );
  AOI220 U74 ( .A(Din[6]), .B(n34), .C(n470), .D(Dout[6]), .Q(n53) );
  AOI220 U75 ( .A(Din[3]), .B(n34), .C(n466), .D(Dout[3]), .Q(n65) );
  AOI220 U76 ( .A(Din[18]), .B(n472), .C(n465), .D(Dout[18]), .Q(n48) );
  AOI220 U77 ( .A(Din[5]), .B(n34), .C(n465), .D(Dout[5]), .Q(n63) );
  AOI220 U78 ( .A(Din[17]), .B(n472), .C(n467), .D(Dout[17]), .Q(n49) );
endmodule


module reg_32 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n303, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491;

  DF3 Dout_reg_31_ ( .D(n460), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n461), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n462), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n463), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n464), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n465), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n466), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n467), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n468), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n469), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n470), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n471), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n472), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n473), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_16_ ( .D(n474), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_15_ ( .D(n475), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n476), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_12_ ( .D(n477), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_11_ ( .D(n478), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_8_ ( .D(n479), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_0_ ( .D(n480), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_7_ ( .D(n481), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_6_ ( .D(n482), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_10_ ( .D(n483), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_13_ ( .D(n485), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_17_ ( .D(n486), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_2_ ( .D(n489), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_3_ ( .D(n491), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_9_ ( .D(n484), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_4_ ( .D(n490), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_5_ ( .D(n487), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_1_ ( .D(n488), .C(Clk), .Q(n303) );
  BUF15 U3 ( .A(n303), .Q(Dout[1]) );
  AOI220 U4 ( .A(Din[25]), .B(n459), .C(n455), .D(Dout[25]), .Q(n41) );
  AOI220 U5 ( .A(Din[24]), .B(n34), .C(n454), .D(Dout[24]), .Q(n42) );
  AOI220 U6 ( .A(Din[23]), .B(n459), .C(n457), .D(Dout[23]), .Q(n43) );
  INV3 U7 ( .A(n458), .Q(n459) );
  CLKBU2 U8 ( .A(n451), .Q(n454) );
  CLKBU2 U9 ( .A(n450), .Q(n452) );
  CLKBU2 U10 ( .A(n450), .Q(n453) );
  CLKBU2 U11 ( .A(n451), .Q(n455) );
  CLKBU2 U12 ( .A(n35), .Q(n456) );
  CLKBU2 U13 ( .A(n35), .Q(n457) );
  INV3 U14 ( .A(n63), .Q(n488) );
  INV3 U15 ( .A(n62), .Q(n487) );
  INV3 U16 ( .A(n66), .Q(n491) );
  INV3 U17 ( .A(n64), .Q(n489) );
  INV3 U18 ( .A(n56), .Q(n481) );
  AOI220 U19 ( .A(Din[7]), .B(n34), .C(n456), .D(Dout[7]), .Q(n56) );
  INV3 U20 ( .A(n52), .Q(n477) );
  AOI220 U21 ( .A(Din[12]), .B(n34), .C(n455), .D(Dout[12]), .Q(n52) );
  INV3 U22 ( .A(n50), .Q(n475) );
  AOI220 U23 ( .A(Din[15]), .B(n34), .C(n453), .D(Dout[15]), .Q(n50) );
  INV3 U24 ( .A(n46), .Q(n471) );
  AOI220 U25 ( .A(Din[20]), .B(n34), .C(n456), .D(Dout[20]), .Q(n46) );
  INV3 U26 ( .A(n44), .Q(n469) );
  AOI220 U27 ( .A(Din[22]), .B(n34), .C(n456), .D(Dout[22]), .Q(n44) );
  INV3 U28 ( .A(n43), .Q(n468) );
  INV3 U29 ( .A(n42), .Q(n467) );
  INV3 U30 ( .A(n57), .Q(n482) );
  AOI220 U31 ( .A(Din[6]), .B(n459), .C(n455), .D(Dout[6]), .Q(n57) );
  INV3 U32 ( .A(n41), .Q(n466) );
  INV3 U33 ( .A(n54), .Q(n479) );
  AOI220 U34 ( .A(Din[8]), .B(n34), .C(n456), .D(Dout[8]), .Q(n54) );
  INV3 U35 ( .A(n40), .Q(n465) );
  AOI221 U36 ( .A(Din[26]), .B(n34), .C(n457), .D(Dout[26]), .Q(n40) );
  INV3 U37 ( .A(n38), .Q(n463) );
  AOI221 U38 ( .A(Din[28]), .B(n34), .C(n453), .D(Dout[28]), .Q(n38) );
  INV3 U39 ( .A(n36), .Q(n461) );
  AOI221 U40 ( .A(Din[30]), .B(n34), .C(n456), .D(Dout[30]), .Q(n36) );
  INV3 U41 ( .A(n61), .Q(n486) );
  AOI220 U42 ( .A(Din[17]), .B(n459), .C(n454), .D(Dout[17]), .Q(n61) );
  INV3 U43 ( .A(n60), .Q(n485) );
  AOI220 U44 ( .A(Din[13]), .B(n34), .C(n454), .D(Dout[13]), .Q(n60) );
  INV3 U45 ( .A(n51), .Q(n476) );
  AOI220 U46 ( .A(Din[14]), .B(n459), .C(n452), .D(Dout[14]), .Q(n51) );
  INV3 U47 ( .A(n49), .Q(n474) );
  AOI220 U48 ( .A(Din[16]), .B(n459), .C(n454), .D(Dout[16]), .Q(n49) );
  INV3 U49 ( .A(n48), .Q(n473) );
  AOI220 U50 ( .A(Din[18]), .B(n34), .C(n452), .D(Dout[18]), .Q(n48) );
  INV3 U51 ( .A(n47), .Q(n472) );
  AOI220 U52 ( .A(Din[19]), .B(n459), .C(n453), .D(Dout[19]), .Q(n47) );
  INV3 U53 ( .A(n45), .Q(n470) );
  AOI220 U54 ( .A(Din[21]), .B(n459), .C(n455), .D(Dout[21]), .Q(n45) );
  INV3 U55 ( .A(n53), .Q(n478) );
  AOI220 U56 ( .A(Din[11]), .B(n459), .C(n457), .D(Dout[11]), .Q(n53) );
  INV3 U57 ( .A(n65), .Q(n490) );
  AOI220 U58 ( .A(Din[4]), .B(n459), .C(n453), .D(Dout[4]), .Q(n65) );
  INV3 U59 ( .A(n59), .Q(n484) );
  AOI220 U60 ( .A(Din[9]), .B(n459), .C(n455), .D(Dout[9]), .Q(n59) );
  INV3 U61 ( .A(n55), .Q(n480) );
  AOI220 U62 ( .A(Din[0]), .B(n459), .C(n457), .D(Dout[0]), .Q(n55) );
  INV3 U63 ( .A(n58), .Q(n483) );
  AOI220 U64 ( .A(Din[10]), .B(n34), .C(n454), .D(Dout[10]), .Q(n58) );
  INV3 U65 ( .A(n39), .Q(n464) );
  AOI221 U66 ( .A(Din[27]), .B(n459), .C(n452), .D(Dout[27]), .Q(n39) );
  INV3 U67 ( .A(n37), .Q(n462) );
  AOI221 U68 ( .A(Din[29]), .B(n459), .C(n454), .D(Dout[29]), .Q(n37) );
  INV3 U69 ( .A(n33), .Q(n460) );
  AOI221 U70 ( .A(Din[31]), .B(n459), .C(n457), .D(Dout[31]), .Q(n33) );
  NOR21 U71 ( .A(Load), .B(Reset), .Q(n450) );
  NOR21 U72 ( .A(Load), .B(Reset), .Q(n451) );
  NOR21 U73 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U74 ( .A(n34), .Q(n458) );
  NOR21 U75 ( .A(n452), .B(Reset), .Q(n34) );
  AOI220 U76 ( .A(Din[1]), .B(n459), .C(n452), .D(Dout[1]), .Q(n63) );
  AOI220 U77 ( .A(Din[5]), .B(n34), .C(n453), .D(Dout[5]), .Q(n62) );
  AOI220 U78 ( .A(Din[2]), .B(n34), .C(n453), .D(Dout[2]), .Q(n64) );
  AOI220 U79 ( .A(Din[3]), .B(n459), .C(n452), .D(Dout[3]), .Q(n66) );
endmodule


module reg_31 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n563, n172, n406, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n511, n512, n513,
         n514, n515, n517, n519, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562;

  DF3 Dout_reg_31_ ( .D(n531), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n532), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n533), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n534), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n535), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n536), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n537), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n538), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n539), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n540), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_3_ ( .D(n544), .C(Clk), .Q(Dout[3]), .QN(n511) );
  DF3 Dout_reg_18_ ( .D(n545), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_19_ ( .D(n546), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_17_ ( .D(n547), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_14_ ( .D(n548), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_21_ ( .D(n549), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_16_ ( .D(n552), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_10_ ( .D(n554), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_8_ ( .D(n555), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_4_ ( .D(n556), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_15_ ( .D(n557), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_13_ ( .D(n558), .C(Clk), .Q(Dout[13]), .QN(n513) );
  DF3 Dout_reg_5_ ( .D(n559), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_9_ ( .D(n562), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_20_ ( .D(n541), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_6_ ( .D(n553), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_2_ ( .D(n560), .C(Clk), .Q(n172) );
  DF3 Dout_reg_7_ ( .D(n542), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_1_ ( .D(n543), .C(Clk), .Q(n406) );
  DF3 Dout_reg_11_ ( .D(n551), .C(Clk), .Q(n563) );
  DF3 Dout_reg_12_ ( .D(n561), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_0_ ( .D(n550), .C(Clk), .Q(Dout[0]) );
  INV8 U3 ( .A(n519), .Q(Dout[11]) );
  INV12 U4 ( .A(n517), .Q(Dout[1]) );
  INV3 U5 ( .A(n511), .Q(n512) );
  INV3 U6 ( .A(n513), .Q(n514) );
  INV6 U7 ( .A(n172), .Q(n515) );
  INV12 U8 ( .A(n515), .Q(Dout[2]) );
  INV6 U9 ( .A(n406), .Q(n517) );
  INV6 U10 ( .A(n563), .Q(n519) );
  AOI220 U11 ( .A(Din[28]), .B(n530), .C(n524), .D(Dout[28]), .Q(n38) );
  AOI220 U12 ( .A(Din[29]), .B(n34), .C(n525), .D(Dout[29]), .Q(n37) );
  INV3 U13 ( .A(n529), .Q(n530) );
  CLKBU2 U14 ( .A(n522), .Q(n525) );
  CLKBU2 U15 ( .A(n521), .Q(n523) );
  CLKBU2 U16 ( .A(n35), .Q(n528) );
  CLKBU2 U17 ( .A(n521), .Q(n524) );
  CLKBU2 U18 ( .A(n522), .Q(n526) );
  CLKBU2 U19 ( .A(n35), .Q(n527) );
  INV3 U20 ( .A(n55), .Q(n551) );
  INV3 U21 ( .A(n47), .Q(n543) );
  INV3 U22 ( .A(n46), .Q(n542) );
  INV3 U23 ( .A(n64), .Q(n560) );
  INV3 U24 ( .A(n57), .Q(n553) );
  INV3 U25 ( .A(n63), .Q(n559) );
  INV3 U26 ( .A(n62), .Q(n558) );
  INV3 U27 ( .A(n59), .Q(n555) );
  INV3 U28 ( .A(n58), .Q(n554) );
  INV3 U29 ( .A(n56), .Q(n552) );
  INV3 U30 ( .A(n51), .Q(n547) );
  INV3 U31 ( .A(n50), .Q(n546) );
  INV3 U32 ( .A(n48), .Q(n544) );
  INV3 U33 ( .A(n65), .Q(n561) );
  AOI220 U34 ( .A(Din[12]), .B(n34), .C(n524), .D(Dout[12]), .Q(n65) );
  INV3 U35 ( .A(n45), .Q(n541) );
  AOI220 U36 ( .A(Din[20]), .B(n34), .C(n526), .D(Dout[20]), .Q(n45) );
  INV3 U37 ( .A(n61), .Q(n557) );
  AOI220 U38 ( .A(Din[15]), .B(n34), .C(n525), .D(Dout[15]), .Q(n61) );
  INV3 U39 ( .A(n53), .Q(n549) );
  AOI220 U40 ( .A(Din[21]), .B(n34), .C(n528), .D(Dout[21]), .Q(n53) );
  INV3 U41 ( .A(n52), .Q(n548) );
  AOI220 U42 ( .A(Din[14]), .B(n530), .C(n526), .D(Dout[14]), .Q(n52) );
  INV3 U43 ( .A(n49), .Q(n545) );
  AOI220 U44 ( .A(Din[18]), .B(n34), .C(n525), .D(Dout[18]), .Q(n49) );
  INV3 U45 ( .A(n44), .Q(n540) );
  AOI220 U46 ( .A(Din[22]), .B(n530), .C(n527), .D(Dout[22]), .Q(n44) );
  INV3 U47 ( .A(n43), .Q(n539) );
  AOI220 U48 ( .A(Din[23]), .B(n34), .C(n528), .D(Dout[23]), .Q(n43) );
  INV3 U49 ( .A(n41), .Q(n537) );
  AOI220 U50 ( .A(Din[25]), .B(n34), .C(n526), .D(Dout[25]), .Q(n41) );
  INV3 U51 ( .A(n39), .Q(n535) );
  AOI220 U52 ( .A(Din[27]), .B(n34), .C(n523), .D(Dout[27]), .Q(n39) );
  INV3 U53 ( .A(n37), .Q(n533) );
  INV3 U54 ( .A(n33), .Q(n531) );
  AOI221 U55 ( .A(Din[31]), .B(n34), .C(n528), .D(Dout[31]), .Q(n33) );
  INV3 U56 ( .A(n66), .Q(n562) );
  AOI220 U57 ( .A(Din[9]), .B(n530), .C(n523), .D(Dout[9]), .Q(n66) );
  INV3 U58 ( .A(n60), .Q(n556) );
  AOI220 U59 ( .A(Din[4]), .B(n530), .C(n525), .D(Dout[4]), .Q(n60) );
  INV3 U60 ( .A(n42), .Q(n538) );
  AOI220 U61 ( .A(Din[24]), .B(n530), .C(n525), .D(Dout[24]), .Q(n42) );
  INV3 U62 ( .A(n40), .Q(n536) );
  AOI220 U63 ( .A(Din[26]), .B(n530), .C(n528), .D(Dout[26]), .Q(n40) );
  INV3 U64 ( .A(n38), .Q(n534) );
  INV3 U65 ( .A(n36), .Q(n532) );
  AOI221 U66 ( .A(Din[30]), .B(n530), .C(n527), .D(Dout[30]), .Q(n36) );
  INV3 U67 ( .A(n54), .Q(n550) );
  AOI220 U68 ( .A(Din[0]), .B(n530), .C(n527), .D(Dout[0]), .Q(n54) );
  NOR21 U69 ( .A(Load), .B(Reset), .Q(n521) );
  NOR21 U70 ( .A(Load), .B(Reset), .Q(n522) );
  NOR21 U71 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U72 ( .A(n34), .Q(n529) );
  NOR21 U73 ( .A(n523), .B(Reset), .Q(n34) );
  AOI220 U74 ( .A(Din[3]), .B(n530), .C(n523), .D(n512), .Q(n48) );
  AOI220 U75 ( .A(Din[10]), .B(n530), .C(n525), .D(Dout[10]), .Q(n58) );
  AOI220 U76 ( .A(Din[19]), .B(n530), .C(n524), .D(Dout[19]), .Q(n50) );
  AOI220 U77 ( .A(Din[8]), .B(n34), .C(n526), .D(Dout[8]), .Q(n59) );
  AOI220 U78 ( .A(Din[2]), .B(n530), .C(n524), .D(Dout[2]), .Q(n64) );
  AOI220 U79 ( .A(Din[1]), .B(n34), .C(n524), .D(Dout[1]), .Q(n47) );
  AOI220 U80 ( .A(Din[16]), .B(n530), .C(n527), .D(Dout[16]), .Q(n56) );
  AOI220 U81 ( .A(Din[13]), .B(n530), .C(n524), .D(n514), .Q(n62) );
  AOI220 U82 ( .A(Din[5]), .B(n34), .C(n523), .D(Dout[5]), .Q(n63) );
  AOI220 U83 ( .A(Din[17]), .B(n34), .C(n523), .D(Dout[17]), .Q(n51) );
  AOI220 U84 ( .A(Din[11]), .B(n34), .C(n528), .D(Dout[11]), .Q(n55) );
  AOI220 U85 ( .A(Din[7]), .B(n530), .C(n527), .D(Dout[7]), .Q(n46) );
  AOI220 U86 ( .A(Din[6]), .B(n530), .C(n526), .D(Dout[6]), .Q(n57) );
endmodule


module reg_30 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n171, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563;

  DF3 Dout_reg_31_ ( .D(n532), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n533), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n534), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n535), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n536), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n537), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n538), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n539), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n540), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n541), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_20_ ( .D(n542), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n543), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_16_ ( .D(n544), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_3_ ( .D(n545), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_8_ ( .D(n546), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_21_ ( .D(n547), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_0_ ( .D(n550), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_11_ ( .D(n551), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_1_ ( .D(n552), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_14_ ( .D(n553), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_5_ ( .D(n554), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_7_ ( .D(n555), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_2_ ( .D(n557), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_12_ ( .D(n558), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_13_ ( .D(n559), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_9_ ( .D(n560), .C(Clk), .Q(n171) );
  DF3 Dout_reg_6_ ( .D(n561), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_17_ ( .D(n562), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_18_ ( .D(n563), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_10_ ( .D(n556), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_15_ ( .D(n549), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_4_ ( .D(n548), .C(Clk), .Q(Dout[4]) );
  CLKBU15 U3 ( .A(n171), .Q(Dout[9]) );
  AOI220 U4 ( .A(Din[28]), .B(n34), .C(n525), .D(Dout[28]), .Q(n38) );
  AOI220 U5 ( .A(Din[29]), .B(n531), .C(n526), .D(Dout[29]), .Q(n37) );
  INV3 U6 ( .A(n530), .Q(n531) );
  CLKBU2 U7 ( .A(n522), .Q(n524) );
  CLKBU2 U8 ( .A(n35), .Q(n529) );
  CLKBU2 U9 ( .A(n522), .Q(n525) );
  CLKBU2 U10 ( .A(n523), .Q(n526) );
  CLKBU2 U11 ( .A(n523), .Q(n527) );
  CLKBU2 U12 ( .A(n35), .Q(n528) );
  INV3 U13 ( .A(n51), .Q(n548) );
  AOI220 U14 ( .A(Din[4]), .B(n531), .C(n524), .D(Dout[4]), .Q(n51) );
  INV3 U15 ( .A(n59), .Q(n556) );
  INV3 U16 ( .A(n65), .Q(n562) );
  INV3 U17 ( .A(n64), .Q(n561) );
  INV3 U18 ( .A(n63), .Q(n560) );
  INV3 U19 ( .A(n62), .Q(n559) );
  INV3 U20 ( .A(n61), .Q(n558) );
  INV3 U21 ( .A(n60), .Q(n557) );
  INV3 U22 ( .A(n58), .Q(n555) );
  INV3 U23 ( .A(n57), .Q(n554) );
  INV3 U24 ( .A(n56), .Q(n553) );
  INV3 U25 ( .A(n55), .Q(n552) );
  INV3 U26 ( .A(n54), .Q(n551) );
  INV3 U27 ( .A(n49), .Q(n546) );
  INV3 U28 ( .A(n48), .Q(n545) );
  INV3 U29 ( .A(n47), .Q(n544) );
  INV3 U30 ( .A(n46), .Q(n543) );
  INV3 U31 ( .A(n66), .Q(n563) );
  AOI220 U32 ( .A(Din[18]), .B(n34), .C(n524), .D(Dout[18]), .Q(n66) );
  INV3 U33 ( .A(n45), .Q(n542) );
  AOI220 U34 ( .A(Din[20]), .B(n531), .C(n527), .D(Dout[20]), .Q(n45) );
  INV3 U35 ( .A(n52), .Q(n549) );
  AOI220 U36 ( .A(Din[15]), .B(n34), .C(n527), .D(Dout[15]), .Q(n52) );
  INV3 U37 ( .A(n53), .Q(n550) );
  AOI220 U38 ( .A(Din[0]), .B(n531), .C(n529), .D(Dout[0]), .Q(n53) );
  INV3 U39 ( .A(n50), .Q(n547) );
  AOI220 U40 ( .A(Din[21]), .B(n34), .C(n525), .D(Dout[21]), .Q(n50) );
  INV3 U41 ( .A(n44), .Q(n541) );
  AOI220 U42 ( .A(Din[22]), .B(n34), .C(n528), .D(Dout[22]), .Q(n44) );
  INV3 U43 ( .A(n43), .Q(n540) );
  AOI220 U44 ( .A(Din[23]), .B(n531), .C(n529), .D(Dout[23]), .Q(n43) );
  INV3 U45 ( .A(n42), .Q(n539) );
  AOI220 U46 ( .A(Din[24]), .B(n34), .C(n526), .D(Dout[24]), .Q(n42) );
  INV3 U47 ( .A(n41), .Q(n538) );
  AOI220 U48 ( .A(Din[25]), .B(n531), .C(n527), .D(Dout[25]), .Q(n41) );
  INV3 U49 ( .A(n40), .Q(n537) );
  AOI220 U50 ( .A(Din[26]), .B(n34), .C(n529), .D(Dout[26]), .Q(n40) );
  INV3 U51 ( .A(n39), .Q(n536) );
  AOI220 U52 ( .A(Din[27]), .B(n531), .C(n524), .D(Dout[27]), .Q(n39) );
  INV3 U53 ( .A(n38), .Q(n535) );
  INV3 U54 ( .A(n37), .Q(n534) );
  INV3 U55 ( .A(n36), .Q(n533) );
  AOI221 U56 ( .A(Din[30]), .B(n34), .C(n528), .D(Dout[30]), .Q(n36) );
  INV3 U57 ( .A(n33), .Q(n532) );
  AOI221 U58 ( .A(Din[31]), .B(n531), .C(n529), .D(Dout[31]), .Q(n33) );
  NOR21 U59 ( .A(Load), .B(Reset), .Q(n522) );
  NOR21 U60 ( .A(Load), .B(Reset), .Q(n523) );
  NOR21 U61 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U62 ( .A(n34), .Q(n530) );
  NOR21 U63 ( .A(n524), .B(Reset), .Q(n34) );
  AOI220 U64 ( .A(Din[3]), .B(n34), .C(n524), .D(Dout[3]), .Q(n48) );
  AOI220 U65 ( .A(Din[10]), .B(n531), .C(n527), .D(Dout[10]), .Q(n59) );
  AOI220 U66 ( .A(Din[12]), .B(n531), .C(n526), .D(Dout[12]), .Q(n61) );
  AOI220 U67 ( .A(Din[19]), .B(n34), .C(n528), .D(Dout[19]), .Q(n46) );
  AOI220 U68 ( .A(Din[8]), .B(n531), .C(n526), .D(Dout[8]), .Q(n49) );
  AOI220 U69 ( .A(Din[14]), .B(n34), .C(n528), .D(Dout[14]), .Q(n56) );
  AOI220 U70 ( .A(Din[16]), .B(n531), .C(n525), .D(Dout[16]), .Q(n47) );
  AOI220 U71 ( .A(Din[5]), .B(n531), .C(n527), .D(Dout[5]), .Q(n57) );
  AOI220 U72 ( .A(Din[9]), .B(n531), .C(n524), .D(Dout[9]), .Q(n63) );
  AOI220 U73 ( .A(Din[2]), .B(n34), .C(n526), .D(Dout[2]), .Q(n60) );
  AOI220 U74 ( .A(Din[17]), .B(n531), .C(n525), .D(Dout[17]), .Q(n65) );
  AOI220 U75 ( .A(Din[11]), .B(n34), .C(n528), .D(Dout[11]), .Q(n54) );
  AOI220 U76 ( .A(Din[7]), .B(n34), .C(n526), .D(Dout[7]), .Q(n58) );
  AOI220 U77 ( .A(Din[1]), .B(n531), .C(n529), .D(Dout[1]), .Q(n55) );
  AOI220 U78 ( .A(Din[13]), .B(n34), .C(n525), .D(Dout[13]), .Q(n62) );
  AOI220 U79 ( .A(Din[6]), .B(n531), .C(n525), .D(Dout[6]), .Q(n64) );
endmodule


module reg_29 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494;

  DF3 Dout_reg_31_ ( .D(n463), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n464), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n465), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n466), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n467), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n468), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n469), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n470), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n471), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n472), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n473), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n474), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n475), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n476), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n477), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_15_ ( .D(n478), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n479), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_13_ ( .D(n480), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_12_ ( .D(n481), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_11_ ( .D(n482), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_10_ ( .D(n483), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_7_ ( .D(n484), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_16_ ( .D(n485), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_0_ ( .D(n486), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_1_ ( .D(n487), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_4_ ( .D(n488), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_6_ ( .D(n490), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_8_ ( .D(n494), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_3_ ( .D(n491), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_2_ ( .D(n489), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_5_ ( .D(n493), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_9_ ( .D(n492), .C(Clk), .Q(Dout[9]) );
  AOI220 U3 ( .A(Din[28]), .B(n34), .C(n456), .D(Dout[28]), .Q(n38) );
  AOI220 U4 ( .A(Din[29]), .B(n462), .C(n457), .D(Dout[29]), .Q(n37) );
  INV3 U5 ( .A(n461), .Q(n462) );
  CLKBU2 U6 ( .A(n453), .Q(n455) );
  CLKBU2 U7 ( .A(n453), .Q(n456) );
  CLKBU2 U8 ( .A(n454), .Q(n457) );
  CLKBU2 U9 ( .A(n35), .Q(n459) );
  CLKBU2 U10 ( .A(n35), .Q(n460) );
  CLKBU2 U11 ( .A(n454), .Q(n458) );
  INV3 U12 ( .A(n63), .Q(n491) );
  AOI220 U13 ( .A(Din[3]), .B(n462), .C(n455), .D(Dout[3]), .Q(n63) );
  INV3 U14 ( .A(n54), .Q(n482) );
  AOI220 U15 ( .A(Din[11]), .B(n34), .C(n459), .D(Dout[11]), .Q(n54) );
  INV3 U16 ( .A(n46), .Q(n474) );
  AOI220 U17 ( .A(Din[20]), .B(n34), .C(n459), .D(Dout[20]), .Q(n46) );
  INV3 U18 ( .A(n57), .Q(n485) );
  AOI220 U19 ( .A(Din[16]), .B(n462), .C(n458), .D(Dout[16]), .Q(n57) );
  INV3 U20 ( .A(n55), .Q(n483) );
  AOI220 U21 ( .A(Din[10]), .B(n462), .C(n460), .D(Dout[10]), .Q(n55) );
  INV3 U22 ( .A(n64), .Q(n492) );
  INV3 U23 ( .A(n65), .Q(n493) );
  INV3 U24 ( .A(n61), .Q(n489) );
  INV3 U25 ( .A(n59), .Q(n487) );
  INV3 U26 ( .A(n53), .Q(n481) );
  INV3 U27 ( .A(n52), .Q(n480) );
  INV3 U28 ( .A(n51), .Q(n479) );
  INV3 U29 ( .A(n49), .Q(n477) );
  INV3 U30 ( .A(n56), .Q(n484) );
  AOI220 U31 ( .A(Din[7]), .B(n34), .C(n459), .D(Dout[7]), .Q(n56) );
  INV3 U32 ( .A(n62), .Q(n490) );
  AOI220 U33 ( .A(Din[6]), .B(n34), .C(n456), .D(Dout[6]), .Q(n62) );
  INV3 U34 ( .A(n58), .Q(n486) );
  AOI220 U35 ( .A(Din[0]), .B(n34), .C(n457), .D(Dout[0]), .Q(n58) );
  INV3 U36 ( .A(n60), .Q(n488) );
  AOI220 U37 ( .A(Din[4]), .B(n34), .C(n457), .D(Dout[4]), .Q(n60) );
  INV3 U38 ( .A(n66), .Q(n494) );
  AOI220 U39 ( .A(Din[8]), .B(n34), .C(n455), .D(Dout[8]), .Q(n66) );
  INV3 U40 ( .A(n50), .Q(n478) );
  AOI220 U41 ( .A(Din[15]), .B(n34), .C(n456), .D(Dout[15]), .Q(n50) );
  INV3 U42 ( .A(n45), .Q(n473) );
  AOI220 U43 ( .A(Din[21]), .B(n462), .C(n458), .D(Dout[21]), .Q(n45) );
  INV3 U44 ( .A(n44), .Q(n472) );
  AOI220 U45 ( .A(Din[22]), .B(n34), .C(n459), .D(Dout[22]), .Q(n44) );
  INV3 U46 ( .A(n42), .Q(n470) );
  AOI220 U47 ( .A(Din[24]), .B(n34), .C(n457), .D(Dout[24]), .Q(n42) );
  INV3 U48 ( .A(n40), .Q(n468) );
  AOI220 U49 ( .A(Din[26]), .B(n34), .C(n460), .D(Dout[26]), .Q(n40) );
  INV3 U50 ( .A(n38), .Q(n466) );
  INV3 U51 ( .A(n36), .Q(n464) );
  AOI221 U52 ( .A(Din[30]), .B(n34), .C(n459), .D(Dout[30]), .Q(n36) );
  INV3 U53 ( .A(n47), .Q(n475) );
  AOI220 U54 ( .A(Din[19]), .B(n462), .C(n456), .D(Dout[19]), .Q(n47) );
  INV3 U55 ( .A(n43), .Q(n471) );
  AOI220 U56 ( .A(Din[23]), .B(n462), .C(n460), .D(Dout[23]), .Q(n43) );
  INV3 U57 ( .A(n41), .Q(n469) );
  AOI220 U58 ( .A(Din[25]), .B(n462), .C(n458), .D(Dout[25]), .Q(n41) );
  INV3 U59 ( .A(n39), .Q(n467) );
  AOI220 U60 ( .A(Din[27]), .B(n462), .C(n455), .D(Dout[27]), .Q(n39) );
  INV3 U61 ( .A(n37), .Q(n465) );
  INV3 U62 ( .A(n33), .Q(n463) );
  AOI221 U63 ( .A(Din[31]), .B(n462), .C(n460), .D(Dout[31]), .Q(n33) );
  INV3 U64 ( .A(n48), .Q(n476) );
  AOI220 U65 ( .A(Din[18]), .B(n34), .C(n455), .D(Dout[18]), .Q(n48) );
  NOR21 U66 ( .A(Load), .B(Reset), .Q(n453) );
  NOR21 U67 ( .A(Load), .B(Reset), .Q(n454) );
  NOR21 U68 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U69 ( .A(n34), .Q(n461) );
  NOR21 U70 ( .A(n455), .B(Reset), .Q(n34) );
  AOI220 U71 ( .A(Din[12]), .B(n462), .C(n460), .D(Dout[12]), .Q(n53) );
  AOI220 U72 ( .A(Din[14]), .B(n462), .C(n455), .D(Dout[14]), .Q(n51) );
  AOI220 U73 ( .A(Din[5]), .B(n462), .C(n456), .D(Dout[5]), .Q(n65) );
  AOI220 U74 ( .A(Din[9]), .B(n34), .C(n456), .D(Dout[9]), .Q(n64) );
  AOI220 U75 ( .A(Din[17]), .B(n462), .C(n457), .D(Dout[17]), .Q(n49) );
  AOI220 U76 ( .A(Din[2]), .B(n462), .C(n457), .D(Dout[2]), .Q(n61) );
  AOI220 U77 ( .A(Din[1]), .B(n462), .C(n458), .D(Dout[1]), .Q(n59) );
  AOI220 U78 ( .A(Din[13]), .B(n462), .C(n458), .D(Dout[13]), .Q(n52) );
endmodule


module reg_28 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n313, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495;

  DF3 Dout_reg_31_ ( .D(n464), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n465), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n466), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n467), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n468), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n469), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n470), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n471), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n472), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n473), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n474), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n475), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n476), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n477), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n478), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_16_ ( .D(n479), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_14_ ( .D(n480), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_13_ ( .D(n481), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_12_ ( .D(n482), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_10_ ( .D(n483), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_9_ ( .D(n484), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_6_ ( .D(n485), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_11_ ( .D(n486), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_0_ ( .D(n487), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_8_ ( .D(n488), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_1_ ( .D(n490), .C(Clk), .Q(Dout[1]), .QN(n450) );
  DF3 Dout_reg_4_ ( .D(n493), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_7_ ( .D(n495), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_15_ ( .D(n492), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_2_ ( .D(n491), .C(Clk), .Q(n313) );
  DF3 Dout_reg_3_ ( .D(n494), .C(Clk), .Q(Dout[3]), .QN(n452) );
  DF3 Dout_reg_5_ ( .D(n489), .C(Clk), .Q(Dout[5]) );
  CLKBU15 U3 ( .A(n313), .Q(Dout[2]) );
  INV3 U4 ( .A(n450), .Q(n451) );
  INV3 U5 ( .A(n452), .Q(n453) );
  AOI220 U6 ( .A(Din[25]), .B(n34), .C(n459), .D(Dout[25]), .Q(n41) );
  AOI220 U7 ( .A(Din[22]), .B(n463), .C(n460), .D(Dout[22]), .Q(n44) );
  AOI220 U8 ( .A(Din[23]), .B(n34), .C(n461), .D(Dout[23]), .Q(n43) );
  AOI220 U9 ( .A(Din[24]), .B(n463), .C(n458), .D(Dout[24]), .Q(n42) );
  INV3 U10 ( .A(n462), .Q(n463) );
  CLKBU2 U11 ( .A(n454), .Q(n456) );
  CLKBU2 U12 ( .A(n454), .Q(n457) );
  CLKBU2 U13 ( .A(n455), .Q(n458) );
  CLKBU2 U14 ( .A(n455), .Q(n459) );
  CLKBU2 U15 ( .A(n35), .Q(n460) );
  CLKBU2 U16 ( .A(n35), .Q(n461) );
  INV3 U17 ( .A(n62), .Q(n491) );
  INV3 U18 ( .A(n66), .Q(n495) );
  INV3 U19 ( .A(n61), .Q(n490) );
  INV3 U20 ( .A(n65), .Q(n494) );
  AOI220 U21 ( .A(Din[3]), .B(n34), .C(n457), .D(n453), .Q(n65) );
  INV3 U22 ( .A(n63), .Q(n492) );
  AOI220 U23 ( .A(Din[15]), .B(n34), .C(n456), .D(Dout[15]), .Q(n63) );
  INV3 U24 ( .A(n59), .Q(n488) );
  AOI220 U25 ( .A(Din[8]), .B(n34), .C(n459), .D(Dout[8]), .Q(n59) );
  INV3 U26 ( .A(n50), .Q(n479) );
  AOI220 U27 ( .A(Din[16]), .B(n463), .C(n457), .D(Dout[16]), .Q(n50) );
  INV3 U28 ( .A(n48), .Q(n477) );
  AOI220 U29 ( .A(Din[18]), .B(n463), .C(n456), .D(Dout[18]), .Q(n48) );
  INV3 U30 ( .A(n47), .Q(n476) );
  AOI220 U31 ( .A(Din[19]), .B(n34), .C(n457), .D(Dout[19]), .Q(n47) );
  INV3 U32 ( .A(n46), .Q(n475) );
  AOI220 U33 ( .A(Din[20]), .B(n463), .C(n460), .D(Dout[20]), .Q(n46) );
  INV3 U34 ( .A(n45), .Q(n474) );
  AOI220 U35 ( .A(Din[21]), .B(n34), .C(n459), .D(Dout[21]), .Q(n45) );
  INV3 U36 ( .A(n44), .Q(n473) );
  INV3 U37 ( .A(n43), .Q(n472) );
  INV3 U38 ( .A(n58), .Q(n487) );
  AOI220 U39 ( .A(Din[0]), .B(n463), .C(n458), .D(Dout[0]), .Q(n58) );
  INV3 U40 ( .A(n42), .Q(n471) );
  INV3 U41 ( .A(n40), .Q(n469) );
  AOI221 U42 ( .A(Din[26]), .B(n463), .C(n461), .D(Dout[26]), .Q(n40) );
  INV3 U43 ( .A(n38), .Q(n467) );
  AOI221 U44 ( .A(Din[28]), .B(n463), .C(n457), .D(Dout[28]), .Q(n38) );
  INV3 U45 ( .A(n36), .Q(n465) );
  AOI221 U46 ( .A(Din[30]), .B(n463), .C(n460), .D(Dout[30]), .Q(n36) );
  INV3 U47 ( .A(n53), .Q(n482) );
  AOI220 U48 ( .A(Din[12]), .B(n34), .C(n461), .D(Dout[12]), .Q(n53) );
  INV3 U49 ( .A(n52), .Q(n481) );
  AOI220 U50 ( .A(Din[13]), .B(n463), .C(n459), .D(Dout[13]), .Q(n52) );
  INV3 U51 ( .A(n51), .Q(n480) );
  AOI220 U52 ( .A(Din[14]), .B(n34), .C(n456), .D(Dout[14]), .Q(n51) );
  INV3 U53 ( .A(n49), .Q(n478) );
  AOI220 U54 ( .A(Din[17]), .B(n34), .C(n458), .D(Dout[17]), .Q(n49) );
  INV3 U55 ( .A(n57), .Q(n486) );
  AOI220 U56 ( .A(Din[11]), .B(n34), .C(n459), .D(Dout[11]), .Q(n57) );
  INV3 U57 ( .A(n64), .Q(n493) );
  AOI220 U58 ( .A(Din[4]), .B(n463), .C(n457), .D(Dout[4]), .Q(n64) );
  INV3 U59 ( .A(n54), .Q(n483) );
  AOI220 U60 ( .A(Din[10]), .B(n463), .C(n460), .D(Dout[10]), .Q(n54) );
  INV3 U61 ( .A(n60), .Q(n489) );
  AOI220 U62 ( .A(Din[5]), .B(n463), .C(n458), .D(Dout[5]), .Q(n60) );
  INV3 U63 ( .A(n55), .Q(n484) );
  AOI220 U64 ( .A(Din[9]), .B(n34), .C(n461), .D(Dout[9]), .Q(n55) );
  INV3 U65 ( .A(n56), .Q(n485) );
  AOI220 U66 ( .A(Din[6]), .B(n463), .C(n460), .D(Dout[6]), .Q(n56) );
  INV3 U67 ( .A(n41), .Q(n470) );
  INV3 U68 ( .A(n39), .Q(n468) );
  AOI221 U69 ( .A(Din[27]), .B(n34), .C(n456), .D(Dout[27]), .Q(n39) );
  INV3 U70 ( .A(n37), .Q(n466) );
  AOI221 U71 ( .A(Din[29]), .B(n34), .C(n458), .D(Dout[29]), .Q(n37) );
  INV3 U72 ( .A(n33), .Q(n464) );
  AOI221 U73 ( .A(Din[31]), .B(n34), .C(n461), .D(Dout[31]), .Q(n33) );
  NOR21 U74 ( .A(Load), .B(Reset), .Q(n454) );
  NOR21 U75 ( .A(Load), .B(Reset), .Q(n455) );
  NOR21 U76 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U77 ( .A(n34), .Q(n462) );
  NOR21 U78 ( .A(n456), .B(Reset), .Q(n34) );
  AOI220 U79 ( .A(Din[1]), .B(n463), .C(n458), .D(n451), .Q(n61) );
  AOI220 U80 ( .A(Din[2]), .B(n463), .C(n457), .D(Dout[2]), .Q(n62) );
  AOI220 U81 ( .A(Din[7]), .B(n463), .C(n456), .D(Dout[7]), .Q(n66) );
endmodule


module reg_27 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n259, n177, n467, n260, n178, n180, n393, n183, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n583, n584, n585, n586, n587, n588, n589, n591, n593, n595,
         n597, n598, n599, n601, n603, n605, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648;

  DF3 Dout_reg_31_ ( .D(n617), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n618), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n619), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n620), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n621), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n622), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n623), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_23_ ( .D(n624), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n625), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n626), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_10_ ( .D(n627), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_24_ ( .D(n629), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_6_ ( .D(n630), .C(Clk), .Q(Dout[6]), .QN(n585) );
  DF3 Dout_reg_3_ ( .D(n632), .C(Clk), .Q(n393) );
  DF3 Dout_reg_12_ ( .D(n633), .C(Clk), .Q(n467) );
  DF3 Dout_reg_9_ ( .D(n634), .C(Clk), .Q(n178) );
  DF3 Dout_reg_15_ ( .D(n635), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_8_ ( .D(n636), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_18_ ( .D(n637), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_7_ ( .D(n638), .C(Clk), .Q(n180) );
  DF3 Dout_reg_20_ ( .D(n640), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_13_ ( .D(n641), .C(Clk), .Q(n177) );
  DF3 Dout_reg_19_ ( .D(n642), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_11_ ( .D(n643), .C(Clk), .Q(n260) );
  DF3 Dout_reg_1_ ( .D(n645), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_16_ ( .D(n646), .C(Clk), .Q(Dout[16]), .QN(n583) );
  DF3 Dout_reg_17_ ( .D(n648), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_4_ ( .D(n647), .C(Clk), .Q(Dout[4]), .QN(n597) );
  DF3 Dout_reg_14_ ( .D(n644), .C(Clk), .Q(n259) );
  DF3 Dout_reg_5_ ( .D(n631), .C(Clk), .Q(Dout[5]), .QN(n587) );
  DF3 Dout_reg_2_ ( .D(n639), .C(Clk), .Q(n183) );
  DF3 Dout_reg_0_ ( .D(n628), .C(Clk), .Q(Dout[0]) );
  INV12 U3 ( .A(n593), .Q(Dout[12]) );
  CLKIN15 U4 ( .A(n601), .Q(Dout[3]) );
  INV12 U5 ( .A(n591), .Q(Dout[11]) );
  CLKIN15 U6 ( .A(n603), .Q(Dout[9]) );
  INV8 U7 ( .A(n595), .Q(Dout[13]) );
  CLKIN12 U8 ( .A(n599), .Q(Dout[2]) );
  INV3 U9 ( .A(n583), .Q(n584) );
  INV3 U10 ( .A(n585), .Q(n586) );
  CLKIN15 U11 ( .A(n605), .Q(Dout[7]) );
  INV3 U12 ( .A(n587), .Q(n588) );
  INV6 U13 ( .A(n180), .Q(n605) );
  CLKIN6 U14 ( .A(n259), .Q(n589) );
  INV12 U15 ( .A(n589), .Q(Dout[14]) );
  CLKIN6 U16 ( .A(n260), .Q(n591) );
  CLKIN6 U17 ( .A(n467), .Q(n593) );
  CLKIN6 U18 ( .A(n177), .Q(n595) );
  INV3 U19 ( .A(n597), .Q(n598) );
  INV6 U20 ( .A(n183), .Q(n599) );
  CLKIN6 U21 ( .A(n393), .Q(n601) );
  CLKIN6 U22 ( .A(n178), .Q(n603) );
  AOI220 U23 ( .A(Din[28]), .B(n616), .C(n610), .D(Dout[28]), .Q(n38) );
  AOI220 U24 ( .A(Din[29]), .B(n34), .C(n611), .D(Dout[29]), .Q(n37) );
  INV3 U25 ( .A(n615), .Q(n616) );
  CLKBU2 U26 ( .A(n608), .Q(n611) );
  CLKBU2 U27 ( .A(n35), .Q(n614) );
  CLKBU2 U28 ( .A(n607), .Q(n609) );
  CLKBU2 U29 ( .A(n607), .Q(n610) );
  CLKBU2 U30 ( .A(n608), .Q(n612) );
  CLKBU2 U31 ( .A(n35), .Q(n613) );
  INV3 U32 ( .A(n57), .Q(n639) );
  INV3 U33 ( .A(n49), .Q(n631) );
  INV3 U34 ( .A(n62), .Q(n644) );
  INV3 U35 ( .A(n65), .Q(n647) );
  INV3 U36 ( .A(n66), .Q(n648) );
  INV3 U37 ( .A(n64), .Q(n646) );
  INV3 U38 ( .A(n63), .Q(n645) );
  INV3 U39 ( .A(n61), .Q(n643) );
  INV3 U40 ( .A(n56), .Q(n638) );
  INV3 U41 ( .A(n54), .Q(n636) );
  INV3 U42 ( .A(n52), .Q(n634) );
  INV3 U43 ( .A(n51), .Q(n633) );
  INV3 U44 ( .A(n50), .Q(n632) );
  INV3 U45 ( .A(n48), .Q(n630) );
  INV3 U46 ( .A(n45), .Q(n627) );
  INV3 U47 ( .A(n44), .Q(n626) );
  INV3 U48 ( .A(n60), .Q(n642) );
  AOI220 U49 ( .A(Din[19]), .B(n616), .C(n611), .D(Dout[19]), .Q(n60) );
  INV3 U50 ( .A(n55), .Q(n637) );
  AOI220 U51 ( .A(Din[18]), .B(n34), .C(n614), .D(Dout[18]), .Q(n55) );
  INV3 U52 ( .A(n47), .Q(n629) );
  AOI220 U53 ( .A(Din[24]), .B(n34), .C(n610), .D(Dout[24]), .Q(n47) );
  INV3 U54 ( .A(n43), .Q(n625) );
  AOI220 U55 ( .A(Din[22]), .B(n34), .C(n614), .D(Dout[22]), .Q(n43) );
  INV3 U56 ( .A(n42), .Q(n624) );
  AOI220 U57 ( .A(Din[23]), .B(n616), .C(n611), .D(Dout[23]), .Q(n42) );
  INV3 U58 ( .A(n41), .Q(n623) );
  AOI220 U59 ( .A(Din[25]), .B(n34), .C(n612), .D(Dout[25]), .Q(n41) );
  INV3 U60 ( .A(n59), .Q(n641) );
  AOI220 U61 ( .A(Din[13]), .B(n34), .C(n612), .D(Dout[13]), .Q(n59) );
  INV3 U62 ( .A(n53), .Q(n635) );
  AOI220 U63 ( .A(Din[15]), .B(n34), .C(n614), .D(Dout[15]), .Q(n53) );
  INV3 U64 ( .A(n39), .Q(n621) );
  AOI220 U65 ( .A(Din[27]), .B(n34), .C(n609), .D(Dout[27]), .Q(n39) );
  INV3 U66 ( .A(n37), .Q(n619) );
  INV3 U67 ( .A(n33), .Q(n617) );
  AOI221 U68 ( .A(Din[31]), .B(n34), .C(n614), .D(Dout[31]), .Q(n33) );
  INV3 U69 ( .A(n46), .Q(n628) );
  AOI220 U70 ( .A(Din[0]), .B(n616), .C(n613), .D(Dout[0]), .Q(n46) );
  INV3 U71 ( .A(n58), .Q(n640) );
  AOI220 U72 ( .A(Din[20]), .B(n616), .C(n611), .D(Dout[20]), .Q(n58) );
  INV3 U73 ( .A(n40), .Q(n622) );
  AOI220 U74 ( .A(Din[26]), .B(n616), .C(n614), .D(Dout[26]), .Q(n40) );
  INV3 U75 ( .A(n38), .Q(n620) );
  INV3 U76 ( .A(n36), .Q(n618) );
  AOI221 U77 ( .A(Din[30]), .B(n616), .C(n613), .D(Dout[30]), .Q(n36) );
  NOR21 U78 ( .A(Load), .B(Reset), .Q(n607) );
  NOR21 U79 ( .A(Load), .B(Reset), .Q(n608) );
  NOR21 U80 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U81 ( .A(n34), .Q(n615) );
  NOR21 U82 ( .A(n609), .B(Reset), .Q(n34) );
  AOI220 U83 ( .A(Din[5]), .B(n34), .C(n611), .D(n588), .Q(n49) );
  AOI220 U84 ( .A(Din[8]), .B(n616), .C(n613), .D(Dout[8]), .Q(n54) );
  AOI220 U85 ( .A(Din[12]), .B(n34), .C(n609), .D(Dout[12]), .Q(n51) );
  AOI220 U86 ( .A(Din[21]), .B(n616), .C(n613), .D(Dout[21]), .Q(n44) );
  AOI220 U87 ( .A(Din[10]), .B(n34), .C(n612), .D(Dout[10]), .Q(n45) );
  AOI220 U88 ( .A(Din[16]), .B(n616), .C(n610), .D(n584), .Q(n64) );
  AOI220 U89 ( .A(Din[1]), .B(n34), .C(n609), .D(Dout[1]), .Q(n63) );
  AOI220 U90 ( .A(Din[11]), .B(n34), .C(n611), .D(Dout[11]), .Q(n61) );
  AOI220 U91 ( .A(Din[3]), .B(n616), .C(n610), .D(Dout[3]), .Q(n50) );
  AOI220 U92 ( .A(Din[7]), .B(n616), .C(n613), .D(Dout[7]), .Q(n56) );
  AOI220 U93 ( .A(Din[17]), .B(n616), .C(n609), .D(Dout[17]), .Q(n66) );
  AOI220 U94 ( .A(Din[6]), .B(n616), .C(n609), .D(n586), .Q(n48) );
  AOI220 U95 ( .A(Din[14]), .B(n616), .C(n610), .D(Dout[14]), .Q(n62) );
  AOI220 U96 ( .A(Din[2]), .B(n34), .C(n612), .D(Dout[2]), .Q(n57) );
  AOI220 U97 ( .A(Din[9]), .B(n616), .C(n612), .D(Dout[9]), .Q(n52) );
  AOI220 U98 ( .A(Din[4]), .B(n616), .C(n610), .D(n598), .Q(n65) );
endmodule


module reg_26 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446;

  DF3 Dout_reg_31_ ( .D(n415), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n416), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n417), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n418), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n419), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n420), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n421), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n422), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n423), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n424), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n425), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n426), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n427), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n428), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n429), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_16_ ( .D(n430), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_15_ ( .D(n431), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n432), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_13_ ( .D(n433), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_12_ ( .D(n434), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_11_ ( .D(n435), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_10_ ( .D(n436), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_9_ ( .D(n437), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_7_ ( .D(n438), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_6_ ( .D(n439), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_5_ ( .D(n440), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_4_ ( .D(n441), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_3_ ( .D(n442), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_2_ ( .D(n443), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_1_ ( .D(n444), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_8_ ( .D(n445), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_0_ ( .D(n446), .C(Clk), .Q(Dout[0]) );
  AOI220 U3 ( .A(Din[28]), .B(n414), .C(n408), .D(Dout[28]), .Q(n38) );
  AOI220 U4 ( .A(Din[29]), .B(n34), .C(n409), .D(Dout[29]), .Q(n37) );
  INV3 U5 ( .A(n413), .Q(n414) );
  CLKBU2 U6 ( .A(n405), .Q(n407) );
  CLKBU2 U7 ( .A(n405), .Q(n408) );
  CLKBU2 U8 ( .A(n35), .Q(n412) );
  CLKBU2 U9 ( .A(n406), .Q(n409) );
  CLKBU2 U10 ( .A(n35), .Q(n411) );
  CLKBU2 U11 ( .A(n406), .Q(n410) );
  INV3 U12 ( .A(n46), .Q(n426) );
  AOI220 U13 ( .A(Din[20]), .B(n414), .C(n411), .D(Dout[20]), .Q(n46) );
  INV3 U14 ( .A(n51), .Q(n431) );
  AOI220 U15 ( .A(Din[15]), .B(n34), .C(n407), .D(Dout[15]), .Q(n51) );
  INV3 U16 ( .A(n47), .Q(n427) );
  AOI220 U17 ( .A(Din[19]), .B(n34), .C(n408), .D(Dout[19]), .Q(n47) );
  INV3 U18 ( .A(n65), .Q(n445) );
  INV3 U19 ( .A(n63), .Q(n443) );
  INV3 U20 ( .A(n62), .Q(n442) );
  INV3 U21 ( .A(n61), .Q(n441) );
  INV3 U22 ( .A(n60), .Q(n440) );
  INV3 U23 ( .A(n59), .Q(n439) );
  INV3 U24 ( .A(n58), .Q(n438) );
  INV3 U25 ( .A(n57), .Q(n437) );
  INV3 U26 ( .A(n56), .Q(n436) );
  INV3 U27 ( .A(n55), .Q(n435) );
  INV3 U28 ( .A(n54), .Q(n434) );
  INV3 U29 ( .A(n52), .Q(n432) );
  INV3 U30 ( .A(n50), .Q(n430) );
  INV3 U31 ( .A(n49), .Q(n429) );
  INV3 U32 ( .A(n45), .Q(n425) );
  INV3 U33 ( .A(n43), .Q(n423) );
  AOI220 U34 ( .A(Din[23]), .B(n34), .C(n412), .D(Dout[23]), .Q(n43) );
  INV3 U35 ( .A(n40), .Q(n420) );
  AOI220 U36 ( .A(Din[26]), .B(n414), .C(n412), .D(Dout[26]), .Q(n40) );
  INV3 U37 ( .A(n39), .Q(n419) );
  AOI220 U38 ( .A(Din[27]), .B(n34), .C(n407), .D(Dout[27]), .Q(n39) );
  INV3 U39 ( .A(n42), .Q(n422) );
  AOI220 U40 ( .A(Din[24]), .B(n414), .C(n409), .D(Dout[24]), .Q(n42) );
  INV3 U41 ( .A(n41), .Q(n421) );
  AOI220 U42 ( .A(Din[25]), .B(n34), .C(n410), .D(Dout[25]), .Q(n41) );
  INV3 U43 ( .A(n66), .Q(n446) );
  AOI220 U44 ( .A(Din[0]), .B(n414), .C(n407), .D(Dout[0]), .Q(n66) );
  INV3 U45 ( .A(n53), .Q(n433) );
  AOI220 U46 ( .A(Din[13]), .B(n34), .C(n412), .D(Dout[13]), .Q(n53) );
  INV3 U47 ( .A(n38), .Q(n418) );
  INV3 U48 ( .A(n64), .Q(n444) );
  AOI220 U49 ( .A(Din[1]), .B(n414), .C(n408), .D(Dout[1]), .Q(n64) );
  INV3 U50 ( .A(n36), .Q(n416) );
  AOI221 U51 ( .A(Din[30]), .B(n414), .C(n411), .D(Dout[30]), .Q(n36) );
  INV3 U52 ( .A(n37), .Q(n417) );
  INV3 U53 ( .A(n33), .Q(n415) );
  AOI221 U54 ( .A(Din[31]), .B(n34), .C(n412), .D(Dout[31]), .Q(n33) );
  INV3 U55 ( .A(n48), .Q(n428) );
  AOI220 U56 ( .A(Din[18]), .B(n414), .C(n407), .D(Dout[18]), .Q(n48) );
  INV3 U57 ( .A(n44), .Q(n424) );
  AOI220 U58 ( .A(Din[22]), .B(n414), .C(n411), .D(Dout[22]), .Q(n44) );
  NOR21 U59 ( .A(Load), .B(Reset), .Q(n405) );
  NOR21 U60 ( .A(Load), .B(Reset), .Q(n406) );
  NOR21 U61 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U62 ( .A(n34), .Q(n413) );
  NOR21 U63 ( .A(n407), .B(Reset), .Q(n34) );
  AOI220 U64 ( .A(Din[5]), .B(n414), .C(n409), .D(Dout[5]), .Q(n60) );
  AOI220 U65 ( .A(Din[8]), .B(n34), .C(n408), .D(Dout[8]), .Q(n65) );
  AOI220 U66 ( .A(Din[12]), .B(n414), .C(n411), .D(Dout[12]), .Q(n54) );
  AOI220 U67 ( .A(Din[21]), .B(n34), .C(n410), .D(Dout[21]), .Q(n45) );
  AOI220 U68 ( .A(Din[10]), .B(n414), .C(n411), .D(Dout[10]), .Q(n56) );
  AOI220 U69 ( .A(Din[16]), .B(n414), .C(n408), .D(Dout[16]), .Q(n50) );
  AOI220 U70 ( .A(Din[11]), .B(n34), .C(n412), .D(Dout[11]), .Q(n55) );
  AOI220 U71 ( .A(Din[7]), .B(n414), .C(n409), .D(Dout[7]), .Q(n58) );
  AOI220 U72 ( .A(Din[3]), .B(n414), .C(n408), .D(Dout[3]), .Q(n62) );
  AOI220 U73 ( .A(Din[17]), .B(n34), .C(n409), .D(Dout[17]), .Q(n49) );
  AOI220 U74 ( .A(Din[6]), .B(n34), .C(n410), .D(Dout[6]), .Q(n59) );
  AOI220 U75 ( .A(Din[14]), .B(n414), .C(n410), .D(Dout[14]), .Q(n52) );
  AOI220 U76 ( .A(Din[2]), .B(n34), .C(n407), .D(Dout[2]), .Q(n63) );
  AOI220 U77 ( .A(Din[9]), .B(n34), .C(n410), .D(Dout[9]), .Q(n57) );
  AOI220 U78 ( .A(Din[4]), .B(n414), .C(n409), .D(Dout[4]), .Q(n61) );
endmodule


module reg_24 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n295, n11, n13, n15, n17, n19, n21, n23, n25, n27, n31, n34, n46, n48,
         n52, n54, n56, n58, n60, n62, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n63,
         n64, n65, n66, n67, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n119, n158, n465, n299, n51, n53,
         n426, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464;

  DF3 Dout_reg_8_ ( .D(n97), .C(Clk), .Q(Dout[8]), .QN(n90) );
  DF3 Dout_reg_7_ ( .D(n98), .C(Clk), .Q(Dout[7]), .QN(n94) );
  DF3 Dout_reg_3_ ( .D(n102), .C(Clk), .Q(Dout[3]), .QN(n92) );
  DF3 Dout_reg_2_ ( .D(n103), .C(Clk), .Q(Dout[2]), .QN(n66) );
  DF3 Dout_reg_0_ ( .D(n105), .C(Clk), .Q(Dout[0]), .QN(n63) );
  DF3 Dout_reg_15_ ( .D(n84), .C(Clk), .Q(Dout[15]), .QN(n19) );
  DF3 Dout_reg_9_ ( .D(n96), .C(Clk), .Q(Dout[9]), .QN(n89) );
  DF3 Dout_reg_4_ ( .D(n101), .C(Clk), .Q(Dout[4]), .QN(n91) );
  DF3 Dout_reg_16_ ( .D(n83), .C(Clk), .Q(Dout[16]), .QN(n21) );
  DF3 Dout_reg_14_ ( .D(n85), .C(Clk), .Q(Dout[14]), .QN(n17) );
  DF3 Dout_reg_6_ ( .D(n99), .C(Clk), .Q(Dout[6]), .QN(n65) );
  DF3 Dout_reg_21_ ( .D(n78), .C(Clk), .Q(Dout[21]), .QN(n31) );
  DF3 Dout_reg_11_ ( .D(n88), .C(Clk), .Q(Dout[11]), .QN(n11) );
  DF3 Dout_reg_1_ ( .D(n104), .C(Clk), .Q(Dout[1]), .QN(n299) );
  DF3 Dout_reg_10_ ( .D(n95), .C(Clk), .Q(n295), .QN(n64) );
  DF3 Dout_reg_13_ ( .D(n86), .C(Clk), .Q(Dout[13]), .QN(n15) );
  DF3 Dout_reg_27_ ( .D(n72), .C(Clk), .Q(Dout[27]), .QN(n54) );
  DF3 Dout_reg_25_ ( .D(n74), .C(Clk), .Q(n465), .QN(n158) );
  DF3 Dout_reg_24_ ( .D(n75), .C(Clk), .Q(Dout[24]), .QN(n48) );
  DF3 Dout_reg_12_ ( .D(n87), .C(Clk), .Q(Dout[12]), .QN(n13) );
  OAI222 U3 ( .A(n65), .B(n429), .C(n431), .D(n458), .Q(n99) );
  OAI222 U4 ( .A(n94), .B(n429), .C(n430), .D(n457), .Q(n98) );
  OAI222 U5 ( .A(n90), .B(n429), .C(n51), .D(n455), .Q(n97) );
  OAI222 U6 ( .A(n89), .B(n429), .C(n431), .D(n456), .Q(n96) );
  OAI222 U7 ( .A(n64), .B(n429), .C(n430), .D(n454), .Q(n95) );
  OAI222 U8 ( .A(n11), .B(n429), .C(n51), .D(n453), .Q(n88) );
  OAI222 U9 ( .A(n429), .B(n13), .C(n431), .D(n452), .Q(n87) );
  OAI222 U10 ( .A(n429), .B(n15), .C(n430), .D(n451), .Q(n86) );
  OAI222 U11 ( .A(n17), .B(n429), .C(n51), .D(n450), .Q(n85) );
  OAI222 U12 ( .A(n19), .B(n429), .C(n431), .D(n449), .Q(n84) );
  OAI222 U13 ( .A(n429), .B(n21), .C(n430), .D(n435), .Q(n83) );
  OAI222 U14 ( .A(n429), .B(n23), .C(n51), .D(n448), .Q(n82) );
  OAI222 U15 ( .A(n25), .B(n429), .C(n431), .D(n433), .Q(n81) );
  OAI222 U16 ( .A(n27), .B(n429), .C(n430), .D(n434), .Q(n80) );
  OAI222 U17 ( .A(n429), .B(n119), .C(n439), .D(n51), .Q(n79) );
  OAI222 U18 ( .A(n31), .B(n429), .C(n431), .D(n438), .Q(n78) );
  OAI222 U19 ( .A(n34), .B(n429), .C(n430), .D(n436), .Q(n77) );
  OAI222 U20 ( .A(n46), .B(n429), .C(n51), .D(n437), .Q(n76) );
  OAI222 U21 ( .A(n48), .B(n429), .C(n440), .D(n431), .Q(n75) );
  OAI222 U22 ( .A(n158), .B(n429), .C(n442), .D(n430), .Q(n74) );
  OAI222 U23 ( .A(n52), .B(n429), .C(n444), .D(n51), .Q(n73) );
  OAI222 U24 ( .A(n54), .B(n429), .C(n431), .D(n441), .Q(n72) );
  OAI222 U25 ( .A(n56), .B(n429), .C(n430), .D(n443), .Q(n71) );
  OAI222 U26 ( .A(n58), .B(n429), .C(n447), .D(n51), .Q(n70) );
  OAI222 U27 ( .A(n60), .B(n429), .C(n431), .D(n446), .Q(n69) );
  OAI222 U28 ( .A(n62), .B(n429), .C(n430), .D(n445), .Q(n68) );
  OAI222 U29 ( .A(n63), .B(n429), .C(n51), .D(n464), .Q(n105) );
  OAI222 U30 ( .A(n299), .B(n429), .C(n431), .D(n463), .Q(n104) );
  OAI222 U31 ( .A(n66), .B(n429), .C(n430), .D(n462), .Q(n103) );
  OAI222 U32 ( .A(n92), .B(n429), .C(n51), .D(n461), .Q(n102) );
  OAI222 U33 ( .A(n91), .B(n429), .C(n431), .D(n460), .Q(n101) );
  OAI222 U34 ( .A(n67), .B(n429), .C(n430), .D(n459), .Q(n100) );
  DF3 Dout_reg_20_ ( .D(n79), .C(Clk), .Q(Dout[20]), .QN(n119) );
  DF3 Dout_reg_28_ ( .D(n71), .C(Clk), .Q(Dout[28]), .QN(n56) );
  DF3 Dout_reg_22_ ( .D(n77), .C(Clk), .Q(Dout[22]), .QN(n34) );
  DF3 Dout_reg_19_ ( .D(n80), .C(Clk), .Q(Dout[19]), .QN(n27) );
  DF3 Dout_reg_23_ ( .D(n76), .C(Clk), .Q(Dout[23]), .QN(n46) );
  DF3 Dout_reg_26_ ( .D(n73), .C(Clk), .Q(Dout[26]), .QN(n52) );
  DF3 Dout_reg_17_ ( .D(n82), .C(Clk), .Q(Dout[17]), .QN(n23) );
  DF3 Dout_reg_5_ ( .D(n100), .C(Clk), .Q(Dout[5]), .QN(n67) );
  DF3 Dout_reg_29_ ( .D(n70), .C(Clk), .Q(Dout[29]), .QN(n58) );
  DF1 Dout_reg_31_ ( .D(n68), .C(Clk), .Q(Dout[31]), .QN(n62) );
  DF1 Dout_reg_30_ ( .D(n69), .C(Clk), .Q(Dout[30]), .QN(n60) );
  DF1 Dout_reg_18_ ( .D(n81), .C(Clk), .Q(Dout[18]), .QN(n25) );
  CLKBU12 U35 ( .A(n465), .Q(Dout[25]) );
  INV3 U36 ( .A(Din[29]), .Q(n447) );
  INV2 U37 ( .A(Din[20]), .Q(n439) );
  INV3 U38 ( .A(Din[17]), .Q(n448) );
  INV3 U39 ( .A(Din[18]), .Q(n433) );
  INV3 U40 ( .A(Din[24]), .Q(n440) );
  INV3 U41 ( .A(Din[28]), .Q(n443) );
  INV3 U42 ( .A(Din[31]), .Q(n445) );
  INV3 U43 ( .A(Din[30]), .Q(n446) );
  INV2 U44 ( .A(Din[16]), .Q(n435) );
  INV2 U45 ( .A(Din[4]), .Q(n460) );
  CLKIN3 U46 ( .A(Din[6]), .Q(n458) );
  CLKIN3 U47 ( .A(Din[5]), .Q(n459) );
  INV2 U48 ( .A(Din[8]), .Q(n455) );
  NAND22 U49 ( .A(n432), .B(n429), .Q(n431) );
  NAND22 U50 ( .A(n432), .B(n429), .Q(n430) );
  NAND22 U51 ( .A(n432), .B(n429), .Q(n51) );
  INV3 U52 ( .A(Reset), .Q(n432) );
  INV3 U53 ( .A(n53), .Q(n429) );
  INV3 U54 ( .A(Din[19]), .Q(n434) );
  INV3 U55 ( .A(Din[22]), .Q(n436) );
  INV3 U56 ( .A(Din[9]), .Q(n456) );
  INV3 U57 ( .A(Din[12]), .Q(n452) );
  INV3 U58 ( .A(Din[13]), .Q(n451) );
  INV3 U59 ( .A(Din[10]), .Q(n454) );
  INV3 U60 ( .A(Din[15]), .Q(n449) );
  INV3 U61 ( .A(Din[7]), .Q(n457) );
  INV3 U62 ( .A(Din[1]), .Q(n463) );
  INV3 U63 ( .A(Din[2]), .Q(n462) );
  INV3 U64 ( .A(Din[23]), .Q(n437) );
  INV3 U65 ( .A(Din[11]), .Q(n453) );
  INV3 U66 ( .A(Din[14]), .Q(n450) );
  CLKIN6 U67 ( .A(n295), .Q(n426) );
  INV3 U68 ( .A(Din[3]), .Q(n461) );
  INV3 U69 ( .A(Din[0]), .Q(n464) );
  NOR20 U70 ( .A(Load), .B(Reset), .Q(n53) );
  INV15 U71 ( .A(n426), .Q(Dout[10]) );
  INV3 U72 ( .A(Din[21]), .Q(n438) );
  INV3 U73 ( .A(Din[25]), .Q(n442) );
  INV3 U74 ( .A(Din[27]), .Q(n441) );
  INV3 U75 ( .A(Din[26]), .Q(n444) );
endmodule


module reg_23 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646;

  DF3 Dout_reg_31_ ( .D(n615), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n616), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n617), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n618), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n619), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n620), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n621), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_21_ ( .D(n622), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n623), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n624), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n625), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n626), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_16_ ( .D(n627), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_8_ ( .D(n628), .C(Clk), .Q(Dout[8]), .QN(n600) );
  DF3 Dout_reg_24_ ( .D(n629), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_13_ ( .D(n630), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_10_ ( .D(n633), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_1_ ( .D(n634), .C(Clk), .Q(Dout[1]), .QN(n594) );
  DF3 Dout_reg_12_ ( .D(n635), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_4_ ( .D(n636), .C(Clk), .Q(Dout[4]), .QN(n590) );
  DF3 Dout_reg_23_ ( .D(n638), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_3_ ( .D(n640), .C(Clk), .Q(Dout[3]), .QN(n598) );
  DF3 Dout_reg_11_ ( .D(n641), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_9_ ( .D(n642), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_0_ ( .D(n643), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_5_ ( .D(n644), .C(Clk), .Q(Dout[5]), .QN(n592) );
  DF3 Dout_reg_2_ ( .D(n637), .C(Clk), .Q(Dout[2]), .QN(n596) );
  DF3 Dout_reg_7_ ( .D(n646), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_15_ ( .D(n631), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n632), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_6_ ( .D(n645), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_22_ ( .D(n639), .C(Clk), .Q(Dout[22]) );
  INV3 U3 ( .A(n590), .Q(n591) );
  INV3 U4 ( .A(n592), .Q(n593) );
  INV3 U5 ( .A(n594), .Q(n595) );
  INV3 U6 ( .A(n596), .Q(n597) );
  INV3 U7 ( .A(n598), .Q(n599) );
  INV3 U8 ( .A(n600), .Q(n601) );
  INV3 U9 ( .A(n613), .Q(n614) );
  INV3 U10 ( .A(n34), .Q(n613) );
  NOR21 U11 ( .A(n605), .B(Reset), .Q(n34) );
  INV3 U12 ( .A(n604), .Q(n605) );
  INV3 U13 ( .A(n608), .Q(n609) );
  INV3 U14 ( .A(n604), .Q(n606) );
  INV3 U15 ( .A(n604), .Q(n607) );
  INV3 U16 ( .A(n608), .Q(n610) );
  INV3 U17 ( .A(n608), .Q(n611) );
  INV3 U18 ( .A(n608), .Q(n612) );
  INV3 U19 ( .A(n59), .Q(n639) );
  INV3 U20 ( .A(n65), .Q(n645) );
  INV3 U21 ( .A(n52), .Q(n632) );
  INV3 U22 ( .A(n51), .Q(n631) );
  INV3 U23 ( .A(n66), .Q(n646) );
  INV3 U24 ( .A(n57), .Q(n637) );
  INV3 U25 ( .A(n64), .Q(n644) );
  INV3 U26 ( .A(n63), .Q(n643) );
  INV3 U27 ( .A(n62), .Q(n642) );
  INV3 U28 ( .A(n61), .Q(n641) );
  INV3 U29 ( .A(n60), .Q(n640) );
  INV3 U30 ( .A(n58), .Q(n638) );
  INV3 U31 ( .A(n56), .Q(n636) );
  INV3 U32 ( .A(n55), .Q(n635) );
  INV3 U33 ( .A(n54), .Q(n634) );
  INV3 U34 ( .A(n53), .Q(n633) );
  INV3 U35 ( .A(n50), .Q(n630) );
  INV3 U36 ( .A(n48), .Q(n628) );
  INV3 U37 ( .A(n47), .Q(n627) );
  INV3 U38 ( .A(n46), .Q(n626) );
  INV3 U39 ( .A(n45), .Q(n625) );
  INV3 U40 ( .A(n44), .Q(n624) );
  INV3 U41 ( .A(n43), .Q(n623) );
  INV3 U42 ( .A(n42), .Q(n622) );
  INV3 U43 ( .A(n40), .Q(n620) );
  INV3 U44 ( .A(n39), .Q(n619) );
  AOI220 U45 ( .A(Din[27]), .B(n34), .C(n35), .D(Dout[27]), .Q(n39) );
  INV3 U46 ( .A(n49), .Q(n629) );
  AOI220 U47 ( .A(Din[24]), .B(n34), .C(n609), .D(Dout[24]), .Q(n49) );
  INV3 U48 ( .A(n37), .Q(n617) );
  AOI220 U49 ( .A(Din[29]), .B(n34), .C(n605), .D(Dout[29]), .Q(n37) );
  INV3 U50 ( .A(n38), .Q(n618) );
  AOI220 U51 ( .A(Din[28]), .B(n614), .C(n602), .D(Dout[28]), .Q(n38) );
  INV3 U52 ( .A(n36), .Q(n616) );
  AOI221 U53 ( .A(Din[30]), .B(n614), .C(n606), .D(Dout[30]), .Q(n36) );
  INV3 U54 ( .A(n33), .Q(n615) );
  AOI221 U55 ( .A(Din[31]), .B(n34), .C(n607), .D(Dout[31]), .Q(n33) );
  INV3 U56 ( .A(n41), .Q(n621) );
  AOI220 U57 ( .A(Din[25]), .B(n34), .C(n35), .D(Dout[25]), .Q(n41) );
  INV3 U58 ( .A(n603), .Q(n608) );
  NOR20 U59 ( .A(Load), .B(Reset), .Q(n603) );
  NOR20 U60 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U61 ( .A(n602), .Q(n604) );
  NOR20 U62 ( .A(Load), .B(Reset), .Q(n602) );
  AOI220 U63 ( .A(Din[21]), .B(n614), .C(n612), .D(Dout[21]), .Q(n42) );
  AOI220 U64 ( .A(Din[20]), .B(n34), .C(n603), .D(Dout[20]), .Q(n43) );
  AOI220 U65 ( .A(Din[26]), .B(n614), .C(n35), .D(Dout[26]), .Q(n40) );
  AOI220 U66 ( .A(Din[19]), .B(n614), .C(n612), .D(Dout[19]), .Q(n44) );
  AOI220 U67 ( .A(Din[18]), .B(n34), .C(n611), .D(Dout[18]), .Q(n45) );
  AOI220 U68 ( .A(Din[12]), .B(n34), .C(n610), .D(Dout[12]), .Q(n55) );
  AOI220 U69 ( .A(Din[14]), .B(n614), .C(n606), .D(Dout[14]), .Q(n52) );
  AOI220 U70 ( .A(Din[13]), .B(n614), .C(n610), .D(Dout[13]), .Q(n50) );
  AOI220 U71 ( .A(Din[4]), .B(n614), .C(n609), .D(n591), .Q(n56) );
  AOI220 U72 ( .A(Din[23]), .B(n614), .C(n606), .D(Dout[23]), .Q(n58) );
  AOI220 U73 ( .A(Din[0]), .B(n34), .C(n611), .D(Dout[0]), .Q(n63) );
  AOI220 U74 ( .A(Din[10]), .B(n34), .C(n605), .D(Dout[10]), .Q(n53) );
  AOI220 U75 ( .A(Din[16]), .B(n34), .C(n611), .D(Dout[16]), .Q(n47) );
  AOI220 U76 ( .A(Din[2]), .B(n34), .C(n611), .D(n597), .Q(n57) );
  AOI220 U77 ( .A(Din[8]), .B(n614), .C(n610), .D(n601), .Q(n48) );
  AOI220 U78 ( .A(Din[5]), .B(n614), .C(n610), .D(n593), .Q(n64) );
  AOI220 U79 ( .A(Din[9]), .B(n614), .C(n612), .D(Dout[9]), .Q(n62) );
  AOI220 U80 ( .A(Din[17]), .B(n614), .C(n607), .D(Dout[17]), .Q(n46) );
  AOI220 U81 ( .A(Din[22]), .B(n34), .C(n609), .D(Dout[22]), .Q(n59) );
  AOI220 U82 ( .A(Din[1]), .B(n614), .C(n35), .D(n595), .Q(n54) );
  AOI220 U83 ( .A(Din[7]), .B(n614), .C(n612), .D(Dout[7]), .Q(n66) );
  AOI220 U84 ( .A(Din[6]), .B(n34), .C(n609), .D(Dout[6]), .Q(n65) );
  AOI220 U85 ( .A(Din[3]), .B(n614), .C(n603), .D(n599), .Q(n60) );
  AOI220 U86 ( .A(Din[11]), .B(n34), .C(n602), .D(Dout[11]), .Q(n61) );
  AOI220 U87 ( .A(Din[15]), .B(n614), .C(n607), .D(Dout[15]), .Q(n51) );
endmodule


module reg_22 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n468, n193, n194, n195, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n582, n584,
         n587, n588, n589, n590, n591, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637;

  DF3 Dout_reg_31_ ( .D(n606), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n607), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n608), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n609), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n610), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n611), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_24_ ( .D(n612), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_21_ ( .D(n613), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n614), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_18_ ( .D(n615), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n616), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_0_ ( .D(n620), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_22_ ( .D(n621), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_23_ ( .D(n622), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_15_ ( .D(n623), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_4_ ( .D(n626), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_2_ ( .D(n627), .C(Clk), .Q(n194) );
  DF3 Dout_reg_12_ ( .D(n629), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_1_ ( .D(n630), .C(Clk), .Q(n195) );
  DF3 Dout_reg_8_ ( .D(n632), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_3_ ( .D(n633), .C(Clk), .Q(n193) );
  DF3 Dout_reg_13_ ( .D(n634), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_19_ ( .D(n635), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_6_ ( .D(n636), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_25_ ( .D(n637), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_16_ ( .D(n617), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_10_ ( .D(n628), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_14_ ( .D(n618), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_11_ ( .D(n624), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_9_ ( .D(n631), .C(Clk), .Q(Dout[9]), .QN(n589) );
  DF3 Dout_reg_7_ ( .D(n625), .C(Clk), .Q(n468) );
  DF3 Dout_reg_5_ ( .D(n619), .C(Clk), .Q(Dout[5]), .QN(n587) );
  CLKBU12 U3 ( .A(n468), .Q(Dout[7]) );
  CLKIN6 U4 ( .A(n194), .Q(n582) );
  INV12 U5 ( .A(n582), .Q(Dout[2]) );
  INV6 U6 ( .A(n195), .Q(n584) );
  INV12 U7 ( .A(n584), .Q(Dout[1]) );
  INV12 U8 ( .A(n591), .Q(Dout[3]) );
  INV3 U9 ( .A(n587), .Q(n588) );
  INV3 U10 ( .A(n589), .Q(n590) );
  CLKIN6 U11 ( .A(n193), .Q(n591) );
  AOI220 U12 ( .A(Din[28]), .B(n605), .C(n601), .D(Dout[28]), .Q(n38) );
  AOI220 U13 ( .A(Din[29]), .B(n34), .C(n596), .D(Dout[29]), .Q(n37) );
  INV3 U14 ( .A(n604), .Q(n605) );
  INV3 U15 ( .A(n34), .Q(n604) );
  NOR21 U16 ( .A(n596), .B(Reset), .Q(n34) );
  INV3 U17 ( .A(n595), .Q(n596) );
  INV3 U18 ( .A(n599), .Q(n600) );
  INV3 U19 ( .A(n595), .Q(n597) );
  INV3 U20 ( .A(n595), .Q(n598) );
  INV3 U21 ( .A(n599), .Q(n601) );
  INV3 U22 ( .A(n599), .Q(n602) );
  INV3 U23 ( .A(n599), .Q(n603) );
  INV3 U24 ( .A(n47), .Q(n618) );
  AOI220 U25 ( .A(Din[14]), .B(n34), .C(n602), .D(Dout[14]), .Q(n47) );
  INV3 U26 ( .A(n65), .Q(n636) );
  AOI220 U27 ( .A(Din[6]), .B(n34), .C(n600), .D(Dout[6]), .Q(n65) );
  INV3 U28 ( .A(n59), .Q(n630) );
  AOI220 U29 ( .A(Din[1]), .B(n34), .C(n593), .D(Dout[1]), .Q(n59) );
  INV3 U30 ( .A(n55), .Q(n626) );
  AOI220 U31 ( .A(Din[4]), .B(n34), .C(n601), .D(Dout[4]), .Q(n55) );
  INV3 U32 ( .A(n49), .Q(n620) );
  AOI220 U33 ( .A(Din[0]), .B(n34), .C(n600), .D(Dout[0]), .Q(n49) );
  INV3 U34 ( .A(n43), .Q(n614) );
  AOI220 U35 ( .A(Din[20]), .B(n34), .C(n35), .D(Dout[20]), .Q(n43) );
  INV3 U36 ( .A(n52), .Q(n623) );
  AOI220 U37 ( .A(Din[15]), .B(n605), .C(n597), .D(Dout[15]), .Q(n52) );
  INV3 U38 ( .A(n44), .Q(n615) );
  AOI220 U39 ( .A(Din[18]), .B(n605), .C(n603), .D(Dout[18]), .Q(n44) );
  INV3 U40 ( .A(n48), .Q(n619) );
  INV3 U41 ( .A(n54), .Q(n625) );
  INV3 U42 ( .A(n60), .Q(n631) );
  INV3 U43 ( .A(n53), .Q(n624) );
  INV3 U44 ( .A(n64), .Q(n635) );
  INV3 U45 ( .A(n63), .Q(n634) );
  INV3 U46 ( .A(n62), .Q(n633) );
  INV3 U47 ( .A(n61), .Q(n632) );
  INV3 U48 ( .A(n58), .Q(n629) );
  INV3 U49 ( .A(n56), .Q(n627) );
  INV3 U50 ( .A(n51), .Q(n622) );
  INV3 U51 ( .A(n50), .Q(n621) );
  INV3 U52 ( .A(n45), .Q(n616) );
  INV3 U53 ( .A(n42), .Q(n613) );
  INV3 U54 ( .A(n66), .Q(n637) );
  AOI220 U55 ( .A(Din[25]), .B(n605), .C(n602), .D(Dout[25]), .Q(n66) );
  INV3 U56 ( .A(n41), .Q(n612) );
  AOI220 U57 ( .A(Din[24]), .B(n34), .C(n594), .D(Dout[24]), .Q(n41) );
  INV3 U58 ( .A(n39), .Q(n610) );
  AOI220 U59 ( .A(Din[27]), .B(n34), .C(n600), .D(Dout[27]), .Q(n39) );
  INV3 U60 ( .A(n38), .Q(n609) );
  INV3 U61 ( .A(n40), .Q(n611) );
  AOI220 U62 ( .A(Din[26]), .B(n605), .C(n35), .D(Dout[26]), .Q(n40) );
  INV3 U63 ( .A(n57), .Q(n628) );
  AOI220 U64 ( .A(Din[10]), .B(n34), .C(n603), .D(Dout[10]), .Q(n57) );
  INV3 U65 ( .A(n46), .Q(n617) );
  AOI220 U66 ( .A(Din[16]), .B(n605), .C(n598), .D(Dout[16]), .Q(n46) );
  INV3 U67 ( .A(n37), .Q(n608) );
  INV3 U68 ( .A(n33), .Q(n606) );
  AOI221 U69 ( .A(Din[31]), .B(n34), .C(n598), .D(Dout[31]), .Q(n33) );
  INV3 U70 ( .A(n36), .Q(n607) );
  AOI221 U71 ( .A(Din[30]), .B(n605), .C(n597), .D(Dout[30]), .Q(n36) );
  INV3 U72 ( .A(n594), .Q(n599) );
  NOR20 U73 ( .A(Load), .B(Reset), .Q(n594) );
  NOR20 U74 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U75 ( .A(n593), .Q(n595) );
  NOR20 U76 ( .A(Load), .B(Reset), .Q(n593) );
  AOI220 U77 ( .A(Din[2]), .B(n605), .C(n600), .D(Dout[2]), .Q(n56) );
  AOI220 U78 ( .A(Din[8]), .B(n34), .C(n593), .D(Dout[8]), .Q(n61) );
  AOI220 U79 ( .A(Din[19]), .B(n605), .C(n601), .D(Dout[19]), .Q(n64) );
  AOI220 U80 ( .A(Din[3]), .B(n605), .C(n603), .D(Dout[3]), .Q(n62) );
  AOI220 U81 ( .A(Din[12]), .B(n605), .C(n597), .D(Dout[12]), .Q(n58) );
  AOI220 U82 ( .A(Din[21]), .B(n605), .C(n603), .D(Dout[21]), .Q(n42) );
  AOI220 U83 ( .A(Din[7]), .B(n605), .C(Dout[7]), .D(n35), .Q(n54) );
  AOI220 U84 ( .A(Din[13]), .B(n34), .C(n602), .D(Dout[13]), .Q(n63) );
  AOI220 U85 ( .A(Din[9]), .B(n605), .C(n594), .D(n590), .Q(n60) );
  AOI220 U86 ( .A(Din[23]), .B(n34), .C(n598), .D(Dout[23]), .Q(n51) );
  AOI220 U87 ( .A(Din[5]), .B(n605), .C(n601), .D(n588), .Q(n48) );
  AOI220 U88 ( .A(Din[17]), .B(n34), .C(n602), .D(Dout[17]), .Q(n45) );
  AOI220 U89 ( .A(Din[22]), .B(n605), .C(n35), .D(Dout[22]), .Q(n50) );
  AOI220 U90 ( .A(Din[11]), .B(n605), .C(n596), .D(Dout[11]), .Q(n53) );
endmodule


module reg_21 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n657, n273, n401, n188, n189, n190, n191, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n593, n595, n597, n598, n599, n600, n601, n602, n603, n605, n607,
         n609, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656;

  DF3 Dout_reg_31_ ( .D(n625), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n626), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n627), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n628), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n629), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n630), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n631), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n632), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n633), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n634), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n635), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_12_ ( .D(n636), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_5_ ( .D(n637), .C(Clk), .Q(n190) );
  DF3 Dout_reg_3_ ( .D(n639), .C(Clk), .Q(n191) );
  DF3 Dout_reg_17_ ( .D(n641), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_7_ ( .D(n642), .C(Clk), .Q(n188) );
  DF3 Dout_reg_15_ ( .D(n643), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_0_ ( .D(n644), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_8_ ( .D(n645), .C(Clk), .Q(Dout[8]), .QN(n597) );
  DF3 Dout_reg_16_ ( .D(n646), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_20_ ( .D(n647), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n649), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_9_ ( .D(n651), .C(Clk), .Q(n401) );
  DF3 Dout_reg_6_ ( .D(n652), .C(Clk), .Q(n189) );
  DF3 Dout_reg_14_ ( .D(n655), .C(Clk), .Q(n657) );
  DF3 Dout_reg_13_ ( .D(n656), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_11_ ( .D(n650), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_2_ ( .D(n654), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_18_ ( .D(n640), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_10_ ( .D(n653), .C(Clk), .Q(n273) );
  DF3 Dout_reg_4_ ( .D(n638), .C(Clk), .Q(Dout[4]), .QN(n601) );
  DF3 Dout_reg_1_ ( .D(n648), .C(Clk), .Q(Dout[1]), .QN(n599) );
  INV12 U3 ( .A(n603), .Q(Dout[10]) );
  CLKBU12 U4 ( .A(n657), .Q(Dout[14]) );
  CLKIN12 U5 ( .A(n595), .Q(Dout[5]) );
  CLKIN15 U6 ( .A(n607), .Q(Dout[7]) );
  INV6 U7 ( .A(n191), .Q(n593) );
  CLKIN15 U8 ( .A(n593), .Q(Dout[3]) );
  INV8 U9 ( .A(n605), .Q(Dout[6]) );
  CLKIN6 U10 ( .A(n190), .Q(n595) );
  INV3 U11 ( .A(n597), .Q(n598) );
  INV3 U12 ( .A(n599), .Q(n600) );
  INV3 U13 ( .A(n601), .Q(n602) );
  INV6 U14 ( .A(n273), .Q(n603) );
  INV6 U15 ( .A(n189), .Q(n605) );
  CLKIN6 U16 ( .A(n188), .Q(n607) );
  CLKIN6 U17 ( .A(n401), .Q(n609) );
  INV12 U18 ( .A(n609), .Q(Dout[9]) );
  AOI220 U19 ( .A(Din[28]), .B(n34), .C(n35), .D(Dout[28]), .Q(n38) );
  AOI220 U20 ( .A(Din[29]), .B(n624), .C(n615), .D(Dout[29]), .Q(n37) );
  INV3 U21 ( .A(n623), .Q(n624) );
  INV3 U22 ( .A(n34), .Q(n623) );
  NOR21 U23 ( .A(n615), .B(Reset), .Q(n34) );
  INV3 U24 ( .A(n614), .Q(n615) );
  INV3 U25 ( .A(n614), .Q(n618) );
  INV3 U26 ( .A(n619), .Q(n622) );
  INV3 U27 ( .A(n619), .Q(n620) );
  INV3 U28 ( .A(n614), .Q(n616) );
  INV3 U29 ( .A(n614), .Q(n617) );
  INV3 U30 ( .A(n619), .Q(n621) );
  INV3 U31 ( .A(n58), .Q(n648) );
  INV3 U32 ( .A(n48), .Q(n638) );
  INV3 U33 ( .A(n63), .Q(n653) );
  INV3 U34 ( .A(n64), .Q(n654) );
  INV3 U35 ( .A(n60), .Q(n650) );
  INV3 U36 ( .A(n66), .Q(n656) );
  INV3 U37 ( .A(n65), .Q(n655) );
  INV3 U38 ( .A(n62), .Q(n652) );
  INV3 U39 ( .A(n61), .Q(n651) );
  INV3 U40 ( .A(n59), .Q(n649) );
  INV3 U41 ( .A(n55), .Q(n645) );
  INV3 U42 ( .A(n54), .Q(n644) );
  INV3 U43 ( .A(n53), .Q(n643) );
  INV3 U44 ( .A(n52), .Q(n642) );
  INV3 U45 ( .A(n51), .Q(n641) );
  INV3 U46 ( .A(n49), .Q(n639) );
  INV3 U47 ( .A(n47), .Q(n637) );
  INV3 U48 ( .A(n46), .Q(n636) );
  INV3 U49 ( .A(n45), .Q(n635) );
  INV3 U50 ( .A(n57), .Q(n647) );
  AOI220 U51 ( .A(Din[20]), .B(n624), .C(n618), .D(Dout[20]), .Q(n57) );
  INV3 U52 ( .A(n50), .Q(n640) );
  AOI220 U53 ( .A(Din[18]), .B(n34), .C(n618), .D(Dout[18]), .Q(n50) );
  INV3 U54 ( .A(n44), .Q(n634) );
  AOI220 U55 ( .A(Din[22]), .B(n34), .C(n622), .D(Dout[22]), .Q(n44) );
  INV3 U56 ( .A(n43), .Q(n633) );
  AOI220 U57 ( .A(Din[23]), .B(n624), .C(n35), .D(Dout[23]), .Q(n43) );
  INV3 U58 ( .A(n42), .Q(n632) );
  AOI220 U59 ( .A(Din[24]), .B(n34), .C(n622), .D(Dout[24]), .Q(n42) );
  INV3 U60 ( .A(n40), .Q(n630) );
  AOI220 U61 ( .A(Din[26]), .B(n34), .C(n35), .D(Dout[26]), .Q(n40) );
  INV3 U62 ( .A(n38), .Q(n628) );
  INV3 U63 ( .A(n36), .Q(n626) );
  AOI221 U64 ( .A(Din[30]), .B(n34), .C(n616), .D(Dout[30]), .Q(n36) );
  INV3 U65 ( .A(n41), .Q(n631) );
  AOI220 U66 ( .A(Din[25]), .B(n624), .C(n613), .D(Dout[25]), .Q(n41) );
  INV3 U67 ( .A(n39), .Q(n629) );
  AOI220 U68 ( .A(Din[27]), .B(n624), .C(n612), .D(Dout[27]), .Q(n39) );
  INV3 U69 ( .A(n37), .Q(n627) );
  INV3 U70 ( .A(n33), .Q(n625) );
  AOI221 U71 ( .A(Din[31]), .B(n624), .C(n617), .D(Dout[31]), .Q(n33) );
  INV3 U72 ( .A(n56), .Q(n646) );
  AOI220 U73 ( .A(Din[16]), .B(n34), .C(n620), .D(Dout[16]), .Q(n56) );
  INV3 U74 ( .A(n613), .Q(n619) );
  NOR20 U75 ( .A(Load), .B(Reset), .Q(n613) );
  NOR20 U76 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U77 ( .A(n612), .Q(n614) );
  NOR20 U78 ( .A(Load), .B(Reset), .Q(n612) );
  AOI220 U79 ( .A(Din[2]), .B(n34), .C(n621), .D(Dout[2]), .Q(n64) );
  AOI220 U80 ( .A(Din[0]), .B(n34), .C(n622), .D(Dout[0]), .Q(n54) );
  AOI220 U81 ( .A(Din[15]), .B(n624), .C(n615), .D(Dout[15]), .Q(n53) );
  AOI220 U82 ( .A(Din[8]), .B(n624), .C(n621), .D(n598), .Q(n55) );
  AOI220 U83 ( .A(Din[19]), .B(n624), .C(n35), .D(Dout[19]), .Q(n59) );
  AOI220 U84 ( .A(Din[12]), .B(n34), .C(n617), .D(Dout[12]), .Q(n46) );
  AOI220 U85 ( .A(Din[21]), .B(n624), .C(n618), .D(Dout[21]), .Q(n45) );
  AOI220 U86 ( .A(Din[6]), .B(n34), .C(n622), .D(Dout[6]), .Q(n62) );
  AOI220 U87 ( .A(Din[7]), .B(n34), .C(n616), .D(Dout[7]), .Q(n52) );
  AOI220 U88 ( .A(Din[4]), .B(n34), .C(n621), .D(n602), .Q(n48) );
  AOI220 U89 ( .A(Din[3]), .B(n624), .C(n620), .D(Dout[3]), .Q(n49) );
  AOI220 U90 ( .A(Din[13]), .B(n34), .C(n618), .D(Dout[13]), .Q(n66) );
  AOI220 U91 ( .A(Din[14]), .B(n624), .C(n620), .D(Dout[14]), .Q(n65) );
  AOI220 U92 ( .A(Din[9]), .B(n624), .C(n612), .D(Dout[9]), .Q(n61) );
  AOI220 U93 ( .A(Din[5]), .B(n624), .C(n620), .D(Dout[5]), .Q(n47) );
  AOI220 U94 ( .A(Din[17]), .B(n624), .C(n617), .D(Dout[17]), .Q(n51) );
  AOI220 U95 ( .A(Din[1]), .B(n34), .C(n616), .D(n600), .Q(n58) );
  AOI220 U96 ( .A(Din[10]), .B(n624), .C(n621), .D(Dout[10]), .Q(n63) );
  AOI220 U97 ( .A(Din[11]), .B(n624), .C(n613), .D(Dout[11]), .Q(n60) );
endmodule


module reg_20 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509;

  DF3 Dout_reg_31_ ( .D(n478), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n479), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n480), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n481), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n482), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n483), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n484), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n485), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_22_ ( .D(n487), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n488), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_19_ ( .D(n489), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_16_ ( .D(n491), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_12_ ( .D(n492), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_10_ ( .D(n493), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_1_ ( .D(n494), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_0_ ( .D(n495), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_5_ ( .D(n496), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_17_ ( .D(n497), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_14_ ( .D(n498), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_20_ ( .D(n499), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_15_ ( .D(n500), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_8_ ( .D(n501), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_6_ ( .D(n503), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_11_ ( .D(n504), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_2_ ( .D(n506), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_13_ ( .D(n507), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_23_ ( .D(n486), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_9_ ( .D(n509), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_4_ ( .D(n505), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_3_ ( .D(n502), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_7_ ( .D(n508), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_18_ ( .D(n490), .C(Clk), .Q(Dout[18]) );
  AOI220 U3 ( .A(Din[27]), .B(n477), .C(n35), .D(Dout[27]), .Q(n39) );
  INV3 U4 ( .A(n476), .Q(n477) );
  INV3 U5 ( .A(n34), .Q(n476) );
  NOR21 U6 ( .A(n468), .B(Reset), .Q(n34) );
  INV3 U7 ( .A(n467), .Q(n468) );
  INV3 U8 ( .A(n471), .Q(n474) );
  INV3 U9 ( .A(n471), .Q(n472) );
  INV3 U10 ( .A(n471), .Q(n475) );
  INV3 U11 ( .A(n467), .Q(n469) );
  INV3 U12 ( .A(n467), .Q(n470) );
  INV3 U13 ( .A(n471), .Q(n473) );
  INV3 U14 ( .A(n48), .Q(n491) );
  AOI220 U15 ( .A(Din[16]), .B(n34), .C(n473), .D(Dout[16]), .Q(n48) );
  INV3 U16 ( .A(n65), .Q(n508) );
  INV3 U17 ( .A(n59), .Q(n502) );
  INV3 U18 ( .A(n62), .Q(n505) );
  INV3 U19 ( .A(n66), .Q(n509) );
  INV3 U20 ( .A(n64), .Q(n507) );
  INV3 U21 ( .A(n61), .Q(n504) );
  INV3 U22 ( .A(n60), .Q(n503) );
  INV3 U23 ( .A(n57), .Q(n500) );
  INV3 U24 ( .A(n55), .Q(n498) );
  INV3 U25 ( .A(n53), .Q(n496) );
  INV3 U26 ( .A(n52), .Q(n495) );
  INV3 U27 ( .A(n51), .Q(n494) );
  INV3 U28 ( .A(n50), .Q(n493) );
  INV3 U29 ( .A(n43), .Q(n486) );
  AOI220 U30 ( .A(Din[23]), .B(n477), .C(n35), .D(Dout[23]), .Q(n43) );
  INV3 U31 ( .A(n56), .Q(n499) );
  AOI220 U32 ( .A(Din[20]), .B(n34), .C(n472), .D(Dout[20]), .Q(n56) );
  INV3 U33 ( .A(n42), .Q(n485) );
  AOI220 U34 ( .A(Din[24]), .B(n34), .C(n475), .D(Dout[24]), .Q(n42) );
  INV3 U35 ( .A(n41), .Q(n484) );
  AOI220 U36 ( .A(Din[25]), .B(n477), .C(n466), .D(Dout[25]), .Q(n41) );
  INV3 U37 ( .A(n54), .Q(n497) );
  AOI220 U38 ( .A(Din[17]), .B(n34), .C(n472), .D(Dout[17]), .Q(n54) );
  INV3 U39 ( .A(n45), .Q(n488) );
  AOI220 U40 ( .A(Din[21]), .B(n477), .C(n474), .D(Dout[21]), .Q(n45) );
  INV3 U41 ( .A(n44), .Q(n487) );
  AOI220 U42 ( .A(Din[22]), .B(n34), .C(n475), .D(Dout[22]), .Q(n44) );
  INV3 U43 ( .A(n47), .Q(n490) );
  AOI220 U44 ( .A(Din[18]), .B(n477), .C(n474), .D(Dout[18]), .Q(n47) );
  INV3 U45 ( .A(n63), .Q(n506) );
  AOI220 U46 ( .A(Din[2]), .B(n477), .C(n474), .D(Dout[2]), .Q(n63) );
  INV3 U47 ( .A(n58), .Q(n501) );
  AOI220 U48 ( .A(Din[8]), .B(n34), .C(n469), .D(Dout[8]), .Q(n58) );
  INV3 U49 ( .A(n40), .Q(n483) );
  AOI220 U50 ( .A(Din[26]), .B(n34), .C(n465), .D(Dout[26]), .Q(n40) );
  INV3 U51 ( .A(n39), .Q(n482) );
  INV3 U52 ( .A(n38), .Q(n481) );
  AOI221 U53 ( .A(Din[28]), .B(n34), .C(n35), .D(Dout[28]), .Q(n38) );
  INV3 U54 ( .A(n46), .Q(n489) );
  AOI220 U55 ( .A(Din[19]), .B(n34), .C(n470), .D(Dout[19]), .Q(n46) );
  INV3 U56 ( .A(n36), .Q(n479) );
  AOI221 U57 ( .A(Din[30]), .B(n34), .C(n469), .D(Dout[30]), .Q(n36) );
  INV3 U58 ( .A(n49), .Q(n492) );
  AOI220 U59 ( .A(Din[12]), .B(n477), .C(n472), .D(Dout[12]), .Q(n49) );
  INV3 U60 ( .A(n37), .Q(n480) );
  AOI221 U61 ( .A(Din[29]), .B(n477), .C(n468), .D(Dout[29]), .Q(n37) );
  INV3 U62 ( .A(n33), .Q(n478) );
  AOI221 U63 ( .A(Din[31]), .B(n477), .C(n470), .D(Dout[31]), .Q(n33) );
  INV3 U64 ( .A(n466), .Q(n471) );
  NOR20 U65 ( .A(Load), .B(Reset), .Q(n466) );
  NOR20 U66 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U67 ( .A(n465), .Q(n467) );
  NOR20 U68 ( .A(Load), .B(Reset), .Q(n465) );
  AOI220 U69 ( .A(Din[0]), .B(n34), .C(n469), .D(Dout[0]), .Q(n52) );
  AOI220 U70 ( .A(Din[15]), .B(n477), .C(n475), .D(Dout[15]), .Q(n57) );
  AOI220 U71 ( .A(Din[11]), .B(n477), .C(n465), .D(Dout[11]), .Q(n61) );
  AOI220 U72 ( .A(Din[9]), .B(n34), .C(n473), .D(Dout[9]), .Q(n66) );
  AOI220 U73 ( .A(Din[7]), .B(n477), .C(n472), .D(Dout[7]), .Q(n65) );
  AOI220 U74 ( .A(Din[5]), .B(n477), .C(n468), .D(Dout[5]), .Q(n53) );
  AOI220 U75 ( .A(Din[6]), .B(n34), .C(n474), .D(Dout[6]), .Q(n60) );
  AOI220 U76 ( .A(Din[4]), .B(n34), .C(n475), .D(Dout[4]), .Q(n62) );
  AOI220 U77 ( .A(Din[13]), .B(n34), .C(n473), .D(Dout[13]), .Q(n64) );
  AOI220 U78 ( .A(Din[3]), .B(n477), .C(n466), .D(Dout[3]), .Q(n59) );
  AOI220 U79 ( .A(Din[14]), .B(n477), .C(n473), .D(Dout[14]), .Q(n55) );
  AOI220 U80 ( .A(Din[1]), .B(n477), .C(n470), .D(Dout[1]), .Q(n51) );
  AOI220 U81 ( .A(Din[10]), .B(n477), .C(n35), .D(Dout[10]), .Q(n50) );
endmodule


module reg_19 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n420, n592, n257, n593, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n532, n533,
         n534, n536, n537, n538, n540, n541, n542, n544, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591;

  DF3 Dout_reg_31_ ( .D(n560), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n561), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n562), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n563), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n564), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n565), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n566), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n567), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n568), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n569), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_20_ ( .D(n570), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_18_ ( .D(n571), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n572), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_16_ ( .D(n573), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_14_ ( .D(n574), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_8_ ( .D(n575), .C(Clk), .Q(n593) );
  DF3 Dout_reg_6_ ( .D(n576), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_2_ ( .D(n577), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_0_ ( .D(n578), .C(Clk), .Q(Dout[0]) );
  DF3 Dout_reg_15_ ( .D(n579), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_7_ ( .D(n580), .C(Clk), .Q(Dout[7]), .QN(n536) );
  DF3 Dout_reg_1_ ( .D(n581), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_21_ ( .D(n582), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_9_ ( .D(n586), .C(Clk), .Q(n257), .QN(n540) );
  DF3 Dout_reg_19_ ( .D(n587), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_3_ ( .D(n590), .C(Clk), .Q(Dout[3]), .QN(n532) );
  DF3 Dout_reg_10_ ( .D(n588), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_4_ ( .D(n591), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_5_ ( .D(n583), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_12_ ( .D(n589), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_11_ ( .D(n584), .C(Clk), .Q(n592) );
  DF3 Dout_reg_13_ ( .D(n585), .C(Clk), .Q(n420) );
  INV8 U3 ( .A(n544), .Q(Dout[9]) );
  INV6 U4 ( .A(n542), .Q(Dout[13]) );
  INV3 U5 ( .A(n420), .Q(n542) );
  CLKIN12 U6 ( .A(n538), .Q(Dout[8]) );
  INV8 U7 ( .A(n534), .Q(Dout[11]) );
  INV3 U8 ( .A(n532), .Q(n533) );
  CLKIN6 U9 ( .A(n592), .Q(n534) );
  INV3 U10 ( .A(n536), .Q(n537) );
  CLKIN6 U11 ( .A(n593), .Q(n538) );
  INV3 U12 ( .A(n540), .Q(n541) );
  CLKIN6 U13 ( .A(n257), .Q(n544) );
  AOI220 U14 ( .A(Din[28]), .B(n558), .C(n546), .D(Dout[28]), .Q(n38) );
  AOI220 U15 ( .A(Din[29]), .B(n559), .C(n549), .D(Dout[29]), .Q(n37) );
  INV3 U16 ( .A(n557), .Q(n558) );
  INV3 U17 ( .A(n557), .Q(n559) );
  INV3 U18 ( .A(n34), .Q(n557) );
  NOR21 U19 ( .A(n549), .B(Reset), .Q(n34) );
  INV3 U20 ( .A(n548), .Q(n549) );
  INV3 U21 ( .A(n553), .Q(n556) );
  INV3 U22 ( .A(n548), .Q(n550) );
  INV3 U23 ( .A(n548), .Q(n551) );
  INV3 U24 ( .A(n548), .Q(n552) );
  INV3 U25 ( .A(n553), .Q(n555) );
  INV3 U26 ( .A(n553), .Q(n554) );
  INV3 U27 ( .A(n60), .Q(n585) );
  INV3 U28 ( .A(n59), .Q(n584) );
  INV3 U29 ( .A(n63), .Q(n588) );
  INV3 U30 ( .A(n56), .Q(n581) );
  INV3 U31 ( .A(n55), .Q(n580) );
  INV3 U32 ( .A(n54), .Q(n579) );
  INV3 U33 ( .A(n49), .Q(n574) );
  INV3 U34 ( .A(n48), .Q(n573) );
  INV3 U35 ( .A(n65), .Q(n590) );
  AOI220 U36 ( .A(Din[3]), .B(n559), .C(n556), .D(n533), .Q(n65) );
  INV3 U37 ( .A(n66), .Q(n591) );
  AOI220 U38 ( .A(Din[4]), .B(n558), .C(n555), .D(Dout[4]), .Q(n66) );
  INV3 U39 ( .A(n62), .Q(n587) );
  AOI220 U40 ( .A(Din[19]), .B(n558), .C(n35), .D(Dout[19]), .Q(n62) );
  INV3 U41 ( .A(n52), .Q(n577) );
  AOI220 U42 ( .A(Din[2]), .B(n558), .C(n551), .D(Dout[2]), .Q(n52) );
  INV3 U43 ( .A(n44), .Q(n569) );
  AOI220 U44 ( .A(Din[22]), .B(n558), .C(n555), .D(Dout[22]), .Q(n44) );
  INV3 U45 ( .A(n41), .Q(n566) );
  AOI220 U46 ( .A(Din[25]), .B(n559), .C(n35), .D(Dout[25]), .Q(n41) );
  INV3 U47 ( .A(n58), .Q(n583) );
  AOI220 U48 ( .A(Din[5]), .B(n558), .C(n550), .D(Dout[5]), .Q(n58) );
  INV3 U49 ( .A(n50), .Q(n575) );
  AOI220 U50 ( .A(Din[8]), .B(n558), .C(n555), .D(Dout[8]), .Q(n50) );
  INV3 U51 ( .A(n47), .Q(n572) );
  AOI220 U52 ( .A(Din[17]), .B(n559), .C(n556), .D(Dout[17]), .Q(n47) );
  INV3 U53 ( .A(n46), .Q(n571) );
  AOI220 U54 ( .A(Din[18]), .B(n558), .C(n554), .D(Dout[18]), .Q(n46) );
  INV3 U55 ( .A(n45), .Q(n570) );
  AOI220 U56 ( .A(Din[20]), .B(n559), .C(n551), .D(Dout[20]), .Q(n45) );
  INV3 U57 ( .A(n43), .Q(n568) );
  AOI220 U58 ( .A(Din[23]), .B(n559), .C(n556), .D(Dout[23]), .Q(n43) );
  INV3 U59 ( .A(n42), .Q(n567) );
  AOI220 U60 ( .A(Din[24]), .B(n558), .C(n547), .D(Dout[24]), .Q(n42) );
  INV3 U61 ( .A(n40), .Q(n565) );
  AOI220 U62 ( .A(Din[26]), .B(n558), .C(n35), .D(Dout[26]), .Q(n40) );
  INV3 U63 ( .A(n39), .Q(n564) );
  AOI220 U64 ( .A(Din[27]), .B(n559), .C(n556), .D(Dout[27]), .Q(n39) );
  INV3 U65 ( .A(n38), .Q(n563) );
  INV3 U66 ( .A(n37), .Q(n562) );
  INV3 U67 ( .A(n36), .Q(n561) );
  AOI221 U68 ( .A(Din[30]), .B(n558), .C(n550), .D(Dout[30]), .Q(n36) );
  INV3 U69 ( .A(n33), .Q(n560) );
  AOI221 U70 ( .A(Din[31]), .B(n559), .C(n551), .D(Dout[31]), .Q(n33) );
  INV3 U71 ( .A(n53), .Q(n578) );
  AOI220 U72 ( .A(Din[0]), .B(n559), .C(n550), .D(Dout[0]), .Q(n53) );
  INV3 U73 ( .A(n51), .Q(n576) );
  AOI220 U74 ( .A(Din[6]), .B(n559), .C(n552), .D(Dout[6]), .Q(n51) );
  INV3 U75 ( .A(n64), .Q(n589) );
  AOI220 U76 ( .A(Din[12]), .B(n558), .C(n546), .D(Dout[12]), .Q(n64) );
  INV3 U77 ( .A(n61), .Q(n586) );
  AOI220 U78 ( .A(Din[9]), .B(n559), .C(n35), .D(n541), .Q(n61) );
  INV3 U79 ( .A(n57), .Q(n582) );
  AOI220 U80 ( .A(Din[21]), .B(n559), .C(n552), .D(Dout[21]), .Q(n57) );
  INV3 U81 ( .A(n547), .Q(n553) );
  NOR20 U82 ( .A(Load), .B(Reset), .Q(n547) );
  NOR20 U83 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U84 ( .A(n546), .Q(n548) );
  NOR20 U85 ( .A(Load), .B(Reset), .Q(n546) );
  AOI220 U86 ( .A(Din[16]), .B(n558), .C(n555), .D(Dout[16]), .Q(n48) );
  AOI220 U87 ( .A(Din[1]), .B(n558), .C(n554), .D(Dout[1]), .Q(n56) );
  AOI220 U88 ( .A(Din[15]), .B(n558), .C(n554), .D(Dout[15]), .Q(n54) );
  AOI220 U89 ( .A(Din[14]), .B(n559), .C(n554), .D(Dout[14]), .Q(n49) );
  AOI220 U90 ( .A(Din[7]), .B(n559), .C(n537), .D(n552), .Q(n55) );
  AOI220 U91 ( .A(Din[10]), .B(n559), .C(n547), .D(Dout[10]), .Q(n63) );
  AOI220 U92 ( .A(Din[11]), .B(n559), .C(n552), .D(Dout[11]), .Q(n59) );
  AOI220 U93 ( .A(Din[13]), .B(n558), .C(n549), .D(Dout[13]), .Q(n60) );
endmodule


module reg_18 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473;

  DF3 Dout_reg_31_ ( .D(n442), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n443), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n444), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n445), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n446), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n447), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n448), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n449), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n450), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n451), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n452), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n453), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n454), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n455), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n456), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_16_ ( .D(n457), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_15_ ( .D(n458), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n459), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_13_ ( .D(n460), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_12_ ( .D(n461), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_11_ ( .D(n462), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_10_ ( .D(n463), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_9_ ( .D(n464), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_8_ ( .D(n465), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_7_ ( .D(n466), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_6_ ( .D(n467), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_5_ ( .D(n468), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_4_ ( .D(n469), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_3_ ( .D(n470), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_2_ ( .D(n471), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_1_ ( .D(n472), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_0_ ( .D(n473), .C(Clk), .Q(Dout[0]) );
  AOI220 U3 ( .A(Din[28]), .B(n34), .C(n429), .D(Dout[28]), .Q(n38) );
  AOI220 U4 ( .A(Din[29]), .B(n441), .C(n432), .D(Dout[29]), .Q(n37) );
  INV3 U5 ( .A(n440), .Q(n441) );
  INV3 U6 ( .A(n34), .Q(n440) );
  NOR21 U7 ( .A(n432), .B(Reset), .Q(n34) );
  INV3 U8 ( .A(n431), .Q(n432) );
  INV3 U9 ( .A(n436), .Q(n438) );
  INV3 U10 ( .A(n436), .Q(n439) );
  INV3 U11 ( .A(n431), .Q(n435) );
  INV3 U12 ( .A(n436), .Q(n437) );
  INV3 U13 ( .A(n431), .Q(n433) );
  INV3 U14 ( .A(n431), .Q(n434) );
  INV3 U15 ( .A(n59), .Q(n466) );
  INV3 U16 ( .A(n56), .Q(n463) );
  INV3 U17 ( .A(n55), .Q(n462) );
  INV3 U18 ( .A(n53), .Q(n460) );
  INV3 U19 ( .A(n52), .Q(n459) );
  INV3 U20 ( .A(n51), .Q(n458) );
  INV3 U21 ( .A(n50), .Q(n457) );
  INV3 U22 ( .A(n66), .Q(n473) );
  AOI220 U23 ( .A(Din[0]), .B(n34), .C(n435), .D(Dout[0]), .Q(n66) );
  INV3 U24 ( .A(n64), .Q(n471) );
  AOI220 U25 ( .A(Din[2]), .B(n34), .C(n435), .D(Dout[2]), .Q(n64) );
  INV3 U26 ( .A(n62), .Q(n469) );
  AOI220 U27 ( .A(Din[4]), .B(n34), .C(n439), .D(Dout[4]), .Q(n62) );
  INV3 U28 ( .A(n60), .Q(n467) );
  AOI220 U29 ( .A(Din[6]), .B(n34), .C(n35), .D(Dout[6]), .Q(n60) );
  INV3 U30 ( .A(n47), .Q(n454) );
  AOI220 U31 ( .A(Din[19]), .B(n441), .C(n438), .D(Dout[19]), .Q(n47) );
  INV3 U32 ( .A(n46), .Q(n453) );
  AOI220 U33 ( .A(Din[20]), .B(n34), .C(n434), .D(Dout[20]), .Q(n46) );
  INV3 U34 ( .A(n45), .Q(n452) );
  AOI220 U35 ( .A(Din[21]), .B(n441), .C(n438), .D(Dout[21]), .Q(n45) );
  INV3 U36 ( .A(n44), .Q(n451) );
  AOI220 U37 ( .A(Din[22]), .B(n34), .C(n439), .D(Dout[22]), .Q(n44) );
  INV3 U38 ( .A(n43), .Q(n450) );
  AOI220 U39 ( .A(Din[23]), .B(n441), .C(n35), .D(Dout[23]), .Q(n43) );
  INV3 U40 ( .A(n42), .Q(n449) );
  AOI220 U41 ( .A(Din[24]), .B(n34), .C(n439), .D(Dout[24]), .Q(n42) );
  INV3 U42 ( .A(n41), .Q(n448) );
  AOI220 U43 ( .A(Din[25]), .B(n441), .C(n430), .D(Dout[25]), .Q(n41) );
  INV3 U44 ( .A(n40), .Q(n447) );
  AOI220 U45 ( .A(Din[26]), .B(n34), .C(n438), .D(Dout[26]), .Q(n40) );
  INV3 U46 ( .A(n39), .Q(n446) );
  AOI220 U47 ( .A(Din[27]), .B(n441), .C(n35), .D(Dout[27]), .Q(n39) );
  INV3 U48 ( .A(n38), .Q(n445) );
  INV3 U49 ( .A(n37), .Q(n444) );
  INV3 U50 ( .A(n58), .Q(n465) );
  AOI220 U51 ( .A(Din[8]), .B(n34), .C(n433), .D(Dout[8]), .Q(n58) );
  INV3 U52 ( .A(n54), .Q(n461) );
  AOI220 U53 ( .A(Din[12]), .B(n34), .C(n35), .D(Dout[12]), .Q(n54) );
  INV3 U54 ( .A(n48), .Q(n455) );
  AOI220 U55 ( .A(Din[18]), .B(n34), .C(n439), .D(Dout[18]), .Q(n48) );
  INV3 U56 ( .A(n36), .Q(n443) );
  AOI221 U57 ( .A(Din[30]), .B(n34), .C(n433), .D(Dout[30]), .Q(n36) );
  INV3 U58 ( .A(n63), .Q(n470) );
  AOI220 U59 ( .A(Din[3]), .B(n441), .C(n438), .D(Dout[3]), .Q(n63) );
  INV3 U60 ( .A(n57), .Q(n464) );
  AOI220 U61 ( .A(Din[9]), .B(n441), .C(n435), .D(Dout[9]), .Q(n57) );
  INV3 U62 ( .A(n49), .Q(n456) );
  AOI220 U63 ( .A(Din[17]), .B(n441), .C(n437), .D(Dout[17]), .Q(n49) );
  INV3 U64 ( .A(n33), .Q(n442) );
  AOI221 U65 ( .A(Din[31]), .B(n441), .C(n434), .D(Dout[31]), .Q(n33) );
  INV3 U66 ( .A(n61), .Q(n468) );
  AOI220 U67 ( .A(Din[5]), .B(n441), .C(n429), .D(Dout[5]), .Q(n61) );
  INV3 U68 ( .A(n65), .Q(n472) );
  AOI220 U69 ( .A(Din[1]), .B(n441), .C(n437), .D(Dout[1]), .Q(n65) );
  INV3 U70 ( .A(n430), .Q(n436) );
  NOR20 U71 ( .A(Load), .B(Reset), .Q(n430) );
  NOR20 U72 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U73 ( .A(n429), .Q(n431) );
  NOR20 U74 ( .A(Load), .B(Reset), .Q(n429) );
  AOI220 U75 ( .A(Din[16]), .B(n34), .C(n435), .D(Dout[16]), .Q(n50) );
  AOI220 U76 ( .A(Din[15]), .B(n441), .C(n434), .D(Dout[15]), .Q(n51) );
  AOI220 U77 ( .A(Din[14]), .B(n34), .C(n433), .D(Dout[14]), .Q(n52) );
  AOI220 U78 ( .A(Din[7]), .B(n441), .C(n430), .D(Dout[7]), .Q(n59) );
  AOI220 U79 ( .A(Din[10]), .B(n441), .C(n437), .D(Dout[10]), .Q(n56) );
  AOI220 U80 ( .A(Din[11]), .B(n441), .C(n437), .D(Dout[11]), .Q(n55) );
  AOI220 U81 ( .A(Din[13]), .B(n441), .C(n432), .D(Dout[13]), .Q(n53) );
endmodule


module reg_17 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437;

  DF3 Dout_reg_31_ ( .D(n406), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n407), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n408), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n409), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n410), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n411), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n412), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n413), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n414), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n415), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n416), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n417), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n418), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n419), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n420), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_16_ ( .D(n421), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_15_ ( .D(n422), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n423), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_13_ ( .D(n424), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_12_ ( .D(n425), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_11_ ( .D(n426), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_10_ ( .D(n427), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_9_ ( .D(n428), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_8_ ( .D(n429), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_7_ ( .D(n430), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_6_ ( .D(n431), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_5_ ( .D(n432), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_4_ ( .D(n433), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_3_ ( .D(n434), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_2_ ( .D(n435), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_1_ ( .D(n436), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_0_ ( .D(n437), .C(Clk), .Q(Dout[0]) );
  INV3 U3 ( .A(n404), .Q(n405) );
  INV3 U4 ( .A(n34), .Q(n404) );
  NOR21 U5 ( .A(n396), .B(Reset), .Q(n34) );
  INV3 U6 ( .A(n395), .Q(n396) );
  INV3 U7 ( .A(n395), .Q(n398) );
  INV3 U8 ( .A(n399), .Q(n400) );
  INV3 U9 ( .A(n399), .Q(n401) );
  INV3 U10 ( .A(n399), .Q(n402) );
  INV3 U11 ( .A(n399), .Q(n403) );
  INV3 U12 ( .A(n395), .Q(n397) );
  INV3 U13 ( .A(n66), .Q(n437) );
  AOI221 U14 ( .A(Din[0]), .B(n405), .C(n398), .D(Dout[0]), .Q(n66) );
  INV3 U15 ( .A(n65), .Q(n436) );
  AOI221 U16 ( .A(Din[1]), .B(n34), .C(n400), .D(Dout[1]), .Q(n65) );
  INV3 U17 ( .A(n64), .Q(n435) );
  AOI221 U18 ( .A(Din[2]), .B(n405), .C(n401), .D(Dout[2]), .Q(n64) );
  INV3 U19 ( .A(n63), .Q(n434) );
  AOI221 U20 ( .A(Din[3]), .B(n34), .C(n402), .D(Dout[3]), .Q(n63) );
  INV3 U21 ( .A(n62), .Q(n433) );
  AOI221 U22 ( .A(Din[4]), .B(n405), .C(n403), .D(Dout[4]), .Q(n62) );
  INV3 U23 ( .A(n61), .Q(n432) );
  AOI221 U24 ( .A(Din[5]), .B(n34), .C(n35), .D(Dout[5]), .Q(n61) );
  INV3 U25 ( .A(n60), .Q(n431) );
  AOI221 U26 ( .A(Din[6]), .B(n405), .C(n394), .D(Dout[6]), .Q(n60) );
  INV3 U27 ( .A(n59), .Q(n430) );
  AOI221 U28 ( .A(Din[7]), .B(n34), .C(n393), .D(Dout[7]), .Q(n59) );
  INV3 U29 ( .A(n58), .Q(n429) );
  AOI221 U30 ( .A(Din[8]), .B(n405), .C(n397), .D(Dout[8]), .Q(n58) );
  INV3 U31 ( .A(n57), .Q(n428) );
  AOI221 U32 ( .A(Din[9]), .B(n34), .C(n398), .D(Dout[9]), .Q(n57) );
  INV3 U33 ( .A(n56), .Q(n427) );
  AOI221 U34 ( .A(Din[10]), .B(n405), .C(n400), .D(Dout[10]), .Q(n56) );
  INV3 U35 ( .A(n55), .Q(n426) );
  AOI221 U36 ( .A(Din[11]), .B(n34), .C(n401), .D(Dout[11]), .Q(n55) );
  INV3 U37 ( .A(n54), .Q(n425) );
  AOI221 U38 ( .A(Din[12]), .B(n405), .C(n35), .D(Dout[12]), .Q(n54) );
  INV3 U39 ( .A(n53), .Q(n424) );
  AOI221 U40 ( .A(Din[13]), .B(n34), .C(n396), .D(Dout[13]), .Q(n53) );
  INV3 U41 ( .A(n52), .Q(n423) );
  AOI221 U42 ( .A(Din[14]), .B(n405), .C(n397), .D(Dout[14]), .Q(n52) );
  INV3 U43 ( .A(n51), .Q(n422) );
  AOI221 U44 ( .A(Din[15]), .B(n34), .C(n401), .D(Dout[15]), .Q(n51) );
  INV3 U45 ( .A(n50), .Q(n421) );
  AOI221 U46 ( .A(Din[16]), .B(n405), .C(n398), .D(Dout[16]), .Q(n50) );
  INV3 U47 ( .A(n49), .Q(n420) );
  AOI221 U48 ( .A(Din[17]), .B(n34), .C(n400), .D(Dout[17]), .Q(n49) );
  INV3 U49 ( .A(n48), .Q(n419) );
  AOI221 U50 ( .A(Din[18]), .B(n405), .C(n401), .D(Dout[18]), .Q(n48) );
  INV3 U51 ( .A(n47), .Q(n418) );
  AOI221 U52 ( .A(Din[19]), .B(n34), .C(n402), .D(Dout[19]), .Q(n47) );
  INV3 U53 ( .A(n46), .Q(n417) );
  AOI221 U54 ( .A(Din[20]), .B(n405), .C(n402), .D(Dout[20]), .Q(n46) );
  INV3 U55 ( .A(n45), .Q(n416) );
  AOI221 U56 ( .A(Din[21]), .B(n34), .C(n402), .D(Dout[21]), .Q(n45) );
  INV3 U57 ( .A(n44), .Q(n415) );
  AOI221 U58 ( .A(Din[22]), .B(n405), .C(n403), .D(Dout[22]), .Q(n44) );
  INV3 U59 ( .A(n43), .Q(n414) );
  AOI221 U60 ( .A(Din[23]), .B(n34), .C(n35), .D(Dout[23]), .Q(n43) );
  INV3 U61 ( .A(n42), .Q(n413) );
  AOI221 U62 ( .A(Din[24]), .B(n405), .C(n403), .D(Dout[24]), .Q(n42) );
  INV3 U63 ( .A(n41), .Q(n412) );
  AOI221 U64 ( .A(Din[25]), .B(n34), .C(n400), .D(Dout[25]), .Q(n41) );
  INV3 U65 ( .A(n40), .Q(n411) );
  AOI221 U66 ( .A(Din[26]), .B(n405), .C(n393), .D(Dout[26]), .Q(n40) );
  INV3 U67 ( .A(n39), .Q(n410) );
  AOI221 U68 ( .A(Din[27]), .B(n34), .C(n35), .D(Dout[27]), .Q(n39) );
  INV3 U69 ( .A(n38), .Q(n409) );
  AOI221 U70 ( .A(Din[28]), .B(n405), .C(n394), .D(Dout[28]), .Q(n38) );
  INV3 U71 ( .A(n37), .Q(n408) );
  AOI221 U72 ( .A(Din[29]), .B(n405), .C(n396), .D(Dout[29]), .Q(n37) );
  INV3 U73 ( .A(n36), .Q(n407) );
  AOI221 U74 ( .A(Din[30]), .B(n405), .C(n397), .D(Dout[30]), .Q(n36) );
  INV3 U75 ( .A(n33), .Q(n406) );
  AOI221 U76 ( .A(Din[31]), .B(n405), .C(n403), .D(Dout[31]), .Q(n33) );
  INV3 U77 ( .A(n394), .Q(n399) );
  NOR20 U78 ( .A(Load), .B(Reset), .Q(n394) );
  NOR20 U79 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U80 ( .A(n393), .Q(n395) );
  NOR20 U81 ( .A(Load), .B(Reset), .Q(n393) );
endmodule


module reg_16 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430;

  DF3 Dout_reg_31_ ( .D(n399), .C(Clk), .Q(Dout[31]) );
  DF3 Dout_reg_30_ ( .D(n400), .C(Clk), .Q(Dout[30]) );
  DF3 Dout_reg_29_ ( .D(n401), .C(Clk), .Q(Dout[29]) );
  DF3 Dout_reg_28_ ( .D(n402), .C(Clk), .Q(Dout[28]) );
  DF3 Dout_reg_27_ ( .D(n403), .C(Clk), .Q(Dout[27]) );
  DF3 Dout_reg_26_ ( .D(n404), .C(Clk), .Q(Dout[26]) );
  DF3 Dout_reg_25_ ( .D(n405), .C(Clk), .Q(Dout[25]) );
  DF3 Dout_reg_24_ ( .D(n406), .C(Clk), .Q(Dout[24]) );
  DF3 Dout_reg_23_ ( .D(n407), .C(Clk), .Q(Dout[23]) );
  DF3 Dout_reg_22_ ( .D(n408), .C(Clk), .Q(Dout[22]) );
  DF3 Dout_reg_21_ ( .D(n409), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_20_ ( .D(n410), .C(Clk), .Q(Dout[20]) );
  DF3 Dout_reg_19_ ( .D(n411), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n412), .C(Clk), .Q(Dout[18]) );
  DF3 Dout_reg_17_ ( .D(n413), .C(Clk), .Q(Dout[17]) );
  DF3 Dout_reg_16_ ( .D(n414), .C(Clk), .Q(Dout[16]) );
  DF3 Dout_reg_15_ ( .D(n415), .C(Clk), .Q(Dout[15]) );
  DF3 Dout_reg_14_ ( .D(n416), .C(Clk), .Q(Dout[14]) );
  DF3 Dout_reg_13_ ( .D(n417), .C(Clk), .Q(Dout[13]) );
  DF3 Dout_reg_12_ ( .D(n418), .C(Clk), .Q(Dout[12]) );
  DF3 Dout_reg_11_ ( .D(n419), .C(Clk), .Q(Dout[11]) );
  DF3 Dout_reg_10_ ( .D(n420), .C(Clk), .Q(Dout[10]) );
  DF3 Dout_reg_9_ ( .D(n421), .C(Clk), .Q(Dout[9]) );
  DF3 Dout_reg_8_ ( .D(n422), .C(Clk), .Q(Dout[8]) );
  DF3 Dout_reg_7_ ( .D(n423), .C(Clk), .Q(Dout[7]) );
  DF3 Dout_reg_6_ ( .D(n424), .C(Clk), .Q(Dout[6]) );
  DF3 Dout_reg_5_ ( .D(n425), .C(Clk), .Q(Dout[5]) );
  DF3 Dout_reg_4_ ( .D(n426), .C(Clk), .Q(Dout[4]) );
  DF3 Dout_reg_3_ ( .D(n427), .C(Clk), .Q(Dout[3]) );
  DF3 Dout_reg_2_ ( .D(n428), .C(Clk), .Q(Dout[2]) );
  DF3 Dout_reg_1_ ( .D(n429), .C(Clk), .Q(Dout[1]) );
  DF3 Dout_reg_0_ ( .D(n430), .C(Clk), .Q(Dout[0]) );
  INV3 U3 ( .A(n397), .Q(n398) );
  INV3 U4 ( .A(n34), .Q(n397) );
  NOR21 U5 ( .A(n389), .B(Reset), .Q(n34) );
  INV3 U6 ( .A(n388), .Q(n389) );
  INV3 U7 ( .A(n388), .Q(n391) );
  INV3 U8 ( .A(n392), .Q(n393) );
  INV3 U9 ( .A(n392), .Q(n394) );
  INV3 U10 ( .A(n392), .Q(n395) );
  INV3 U11 ( .A(n392), .Q(n396) );
  INV3 U12 ( .A(n388), .Q(n390) );
  INV3 U13 ( .A(n66), .Q(n430) );
  AOI221 U14 ( .A(Din[0]), .B(n398), .C(n391), .D(Dout[0]), .Q(n66) );
  INV3 U15 ( .A(n65), .Q(n429) );
  AOI221 U16 ( .A(Din[1]), .B(n34), .C(n393), .D(Dout[1]), .Q(n65) );
  INV3 U17 ( .A(n64), .Q(n428) );
  AOI221 U18 ( .A(Din[2]), .B(n398), .C(n394), .D(Dout[2]), .Q(n64) );
  INV3 U19 ( .A(n63), .Q(n427) );
  AOI221 U20 ( .A(Din[3]), .B(n34), .C(n395), .D(Dout[3]), .Q(n63) );
  INV3 U21 ( .A(n62), .Q(n426) );
  AOI221 U22 ( .A(Din[4]), .B(n398), .C(n396), .D(Dout[4]), .Q(n62) );
  INV3 U23 ( .A(n61), .Q(n425) );
  AOI221 U24 ( .A(Din[5]), .B(n34), .C(n35), .D(Dout[5]), .Q(n61) );
  INV3 U25 ( .A(n60), .Q(n424) );
  AOI221 U26 ( .A(Din[6]), .B(n398), .C(n387), .D(Dout[6]), .Q(n60) );
  INV3 U27 ( .A(n59), .Q(n423) );
  AOI221 U28 ( .A(Din[7]), .B(n34), .C(n386), .D(Dout[7]), .Q(n59) );
  INV3 U29 ( .A(n58), .Q(n422) );
  AOI221 U30 ( .A(Din[8]), .B(n398), .C(n390), .D(Dout[8]), .Q(n58) );
  INV3 U31 ( .A(n57), .Q(n421) );
  AOI221 U32 ( .A(Din[9]), .B(n34), .C(n391), .D(Dout[9]), .Q(n57) );
  INV3 U33 ( .A(n56), .Q(n420) );
  AOI221 U34 ( .A(Din[10]), .B(n398), .C(n393), .D(Dout[10]), .Q(n56) );
  INV3 U35 ( .A(n55), .Q(n419) );
  AOI221 U36 ( .A(Din[11]), .B(n34), .C(n394), .D(Dout[11]), .Q(n55) );
  INV3 U37 ( .A(n54), .Q(n418) );
  AOI221 U38 ( .A(Din[12]), .B(n398), .C(n35), .D(Dout[12]), .Q(n54) );
  INV3 U39 ( .A(n53), .Q(n417) );
  AOI221 U40 ( .A(Din[13]), .B(n34), .C(n389), .D(Dout[13]), .Q(n53) );
  INV3 U41 ( .A(n52), .Q(n416) );
  AOI221 U42 ( .A(Din[14]), .B(n398), .C(n390), .D(Dout[14]), .Q(n52) );
  INV3 U43 ( .A(n51), .Q(n415) );
  AOI221 U44 ( .A(Din[15]), .B(n34), .C(n394), .D(Dout[15]), .Q(n51) );
  INV3 U45 ( .A(n50), .Q(n414) );
  AOI221 U46 ( .A(Din[16]), .B(n398), .C(n391), .D(Dout[16]), .Q(n50) );
  INV3 U47 ( .A(n49), .Q(n413) );
  AOI221 U48 ( .A(Din[17]), .B(n34), .C(n393), .D(Dout[17]), .Q(n49) );
  INV3 U49 ( .A(n48), .Q(n412) );
  AOI221 U50 ( .A(Din[18]), .B(n398), .C(n394), .D(Dout[18]), .Q(n48) );
  INV3 U51 ( .A(n47), .Q(n411) );
  AOI221 U52 ( .A(Din[19]), .B(n34), .C(n395), .D(Dout[19]), .Q(n47) );
  INV3 U53 ( .A(n46), .Q(n410) );
  AOI221 U54 ( .A(Din[20]), .B(n398), .C(n395), .D(Dout[20]), .Q(n46) );
  INV3 U55 ( .A(n45), .Q(n409) );
  AOI221 U56 ( .A(Din[21]), .B(n34), .C(n395), .D(Dout[21]), .Q(n45) );
  INV3 U57 ( .A(n44), .Q(n408) );
  AOI221 U58 ( .A(Din[22]), .B(n398), .C(n396), .D(Dout[22]), .Q(n44) );
  INV3 U59 ( .A(n43), .Q(n407) );
  AOI221 U60 ( .A(Din[23]), .B(n34), .C(n35), .D(Dout[23]), .Q(n43) );
  INV3 U61 ( .A(n42), .Q(n406) );
  AOI221 U62 ( .A(Din[24]), .B(n398), .C(n396), .D(Dout[24]), .Q(n42) );
  INV3 U63 ( .A(n41), .Q(n405) );
  AOI221 U64 ( .A(Din[25]), .B(n34), .C(n393), .D(Dout[25]), .Q(n41) );
  INV3 U65 ( .A(n40), .Q(n404) );
  AOI221 U66 ( .A(Din[26]), .B(n398), .C(n386), .D(Dout[26]), .Q(n40) );
  INV3 U67 ( .A(n39), .Q(n403) );
  AOI221 U68 ( .A(Din[27]), .B(n34), .C(n35), .D(Dout[27]), .Q(n39) );
  INV3 U69 ( .A(n38), .Q(n402) );
  AOI221 U70 ( .A(Din[28]), .B(n398), .C(n387), .D(Dout[28]), .Q(n38) );
  INV3 U71 ( .A(n37), .Q(n401) );
  AOI221 U72 ( .A(Din[29]), .B(n398), .C(n389), .D(Dout[29]), .Q(n37) );
  INV3 U73 ( .A(n36), .Q(n400) );
  AOI221 U74 ( .A(Din[30]), .B(n398), .C(n390), .D(Dout[30]), .Q(n36) );
  INV3 U75 ( .A(n33), .Q(n399) );
  AOI221 U76 ( .A(Din[31]), .B(n398), .C(n396), .D(Dout[31]), .Q(n33) );
  INV3 U77 ( .A(n387), .Q(n392) );
  NOR20 U78 ( .A(Load), .B(Reset), .Q(n387) );
  NOR20 U79 ( .A(Load), .B(Reset), .Q(n35) );
  INV3 U80 ( .A(n386), .Q(n388) );
  NOR20 U81 ( .A(Load), .B(Reset), .Q(n386) );
endmodule


module adder_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n418, n427,
         n436, n437, n443, n444, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n594, n595, n596;

  OAI212 U11 ( .A(n42), .B(n527), .C(n43), .Q(n41) );
  OAI212 U25 ( .A(n53), .B(n527), .C(n54), .Q(n52) );
  OAI212 U51 ( .A(n527), .B(n73), .C(n74), .Q(n72) );
  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U77 ( .A(n91), .B(n527), .C(n92), .Q(n90) );
  OAI212 U91 ( .A(n102), .B(n527), .C(n103), .Q(n101) );
  OAI212 U101 ( .A(n536), .B(n527), .C(n530), .Q(n108) );
  OAI212 U115 ( .A(n120), .B(n527), .C(n121), .Q(n119) );
  OAI212 U127 ( .A(n527), .B(n129), .C(n130), .Q(n128) );
  OAI212 U135 ( .A(n137), .B(n145), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n527), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n527), .B(n158), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n534), .B(n527), .C(n528), .Q(n164) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U207 ( .A(n188), .B(n583), .C(n189), .Q(n187) );
  OAI212 U219 ( .A(n197), .B(n583), .C(n198), .Q(n196) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n583), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n579), .B(n583), .C(n580), .Q(n232) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  AOI212 U321 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U447 ( .A(n274), .B(n591), .C(n275), .Q(n273) );
  AOI212 U387 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U393 ( .A(n5), .B(n514), .C(n71), .Q(n67) );
  OAI222 U398 ( .A(n173), .B(n177), .C(n596), .D(n537), .Q(n172) );
  OAI222 U400 ( .A(n155), .B(n163), .C(n595), .D(n541), .Q(n154) );
  NOR24 U428 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR24 U432 ( .A(n185), .B(n194), .Q(n183) );
  NOR24 U438 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NOR24 U451 ( .A(A[23]), .B(B[23]), .Q(n117) );
  OAI212 U459 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  NOR24 U463 ( .A(A[26]), .B(B[26]), .Q(n88) );
  OAI212 U469 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NOR24 U470 ( .A(A[29]), .B(B[29]), .Q(n61) );
  NOR24 U478 ( .A(A[11]), .B(B[11]), .Q(n223) );
  OAI212 U482 ( .A(n117), .B(n127), .C(n118), .Q(n116) );
  NOR24 U485 ( .A(A[19]), .B(B[19]), .Q(n155) );
  NOR24 U493 ( .A(A[17]), .B(B[17]), .Q(n173) );
  OAI212 U507 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U513 ( .A(n82), .B(n527), .C(n83), .Q(n81) );
  XNR22 U520 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR22 U531 ( .A(n10), .B(n72), .Q(SUM[28]) );
  AOI212 U535 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR24 U539 ( .A(B[22]), .B(A[22]), .Q(n126) );
  OAI212 U431 ( .A(n194), .B(n570), .C(n195), .Q(n191) );
  OAI212 U504 ( .A(n427), .B(n46), .C(n47), .Q(n45) );
  NOR24 U511 ( .A(B[14]), .B(A[14]), .Q(n194) );
  XNR22 U349 ( .A(n26), .B(n214), .Q(SUM[12]) );
  INV6 U350 ( .A(n59), .Q(n560) );
  XNR22 U351 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NOR24 U352 ( .A(A[13]), .B(B[13]), .Q(n205) );
  INV4 U353 ( .A(n247), .Q(n583) );
  XNR22 U354 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND21 U355 ( .A(A[13]), .B(B[13]), .Q(n206) );
  INV0 U356 ( .A(n204), .Q(n570) );
  INV2 U357 ( .A(n573), .Q(n509) );
  INV1 U358 ( .A(n203), .Q(n510) );
  INV3 U359 ( .A(n510), .Q(n511) );
  NOR22 U360 ( .A(A[12]), .B(B[12]), .Q(n212) );
  NAND20 U361 ( .A(n578), .B(n245), .Q(n30) );
  OAI211 U362 ( .A(n208), .B(n583), .C(n209), .Q(n207) );
  XNR22 U363 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND23 U364 ( .A(n239), .B(n221), .Q(n219) );
  NOR23 U365 ( .A(n241), .B(n244), .Q(n239) );
  NAND28 U366 ( .A(n59), .B(n556), .Q(n46) );
  INV8 U367 ( .A(n50), .Q(n556) );
  BUF15 U368 ( .A(n178), .Q(n527) );
  NOR24 U369 ( .A(n162), .B(n155), .Q(n153) );
  NAND26 U370 ( .A(n203), .B(n183), .Q(n181) );
  NOR23 U371 ( .A(n117), .B(n126), .Q(n115) );
  NOR23 U372 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NOR23 U373 ( .A(A[18]), .B(B[18]), .Q(n162) );
  NAND22 U374 ( .A(B[12]), .B(A[12]), .Q(n213) );
  NOR23 U375 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND24 U376 ( .A(n115), .B(n135), .Q(n113) );
  NAND23 U377 ( .A(B[18]), .B(A[18]), .Q(n163) );
  NOR22 U378 ( .A(n173), .B(n176), .Q(n171) );
  NOR23 U379 ( .A(A[7]), .B(B[7]), .Q(n252) );
  NOR23 U380 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND22 U381 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NOR23 U382 ( .A(A[25]), .B(B[25]), .Q(n99) );
  INV3 U383 ( .A(n98), .Q(n550) );
  NAND22 U384 ( .A(B[23]), .B(A[23]), .Q(n118) );
  NAND22 U385 ( .A(B[22]), .B(A[22]), .Q(n127) );
  NOR23 U386 ( .A(n181), .B(n219), .Q(n179) );
  NOR22 U388 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NAND22 U389 ( .A(B[8]), .B(A[8]), .Q(n245) );
  AOI211 U390 ( .A(n589), .B(n258), .C(n259), .Q(n257) );
  NOR22 U391 ( .A(A[6]), .B(B[6]), .Q(n255) );
  NOR22 U392 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U394 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NOR23 U395 ( .A(A[21]), .B(B[21]), .Q(n520) );
  NOR23 U396 ( .A(A[21]), .B(B[21]), .Q(n137) );
  NOR23 U397 ( .A(n113), .B(n151), .Q(n111) );
  NAND23 U399 ( .A(n171), .B(n153), .Q(n151) );
  INV3 U401 ( .A(B[19]), .Q(n595) );
  NOR23 U402 ( .A(A[27]), .B(B[27]), .Q(n79) );
  INV3 U403 ( .A(A[19]), .Q(n541) );
  XOR21 U404 ( .A(n22), .B(n527), .Q(SUM[16]) );
  NAND21 U405 ( .A(n582), .B(n253), .Q(n31) );
  CLKIN0 U406 ( .A(n529), .Q(n522) );
  AOI211 U407 ( .A(n529), .B(n549), .C(n548), .Q(n141) );
  CLKIN0 U408 ( .A(n418), .Q(n528) );
  CLKBU2 U409 ( .A(n240), .Q(n512) );
  NOR24 U410 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND23 U411 ( .A(A[20]), .B(B[20]), .Q(n145) );
  INV3 U412 ( .A(n151), .Q(n535) );
  INV2 U413 ( .A(n136), .Q(n543) );
  AOI212 U414 ( .A(n523), .B(n552), .C(n518), .Q(n103) );
  CLKIN3 U415 ( .A(n163), .Q(n539) );
  BUF2 U416 ( .A(n145), .Q(n513) );
  BUF6 U417 ( .A(n70), .Q(n514) );
  NOR23 U418 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NAND23 U419 ( .A(A[28]), .B(B[28]), .Q(n71) );
  INV3 U420 ( .A(n572), .Q(n515) );
  NAND23 U421 ( .A(n111), .B(n44), .Q(n42) );
  CLKIN3 U422 ( .A(n268), .Q(n589) );
  BUF2 U423 ( .A(n155), .Q(n516) );
  NAND28 U424 ( .A(n526), .B(n80), .Q(n78) );
  NOR23 U425 ( .A(B[24]), .B(A[24]), .Q(n106) );
  INV3 U426 ( .A(n135), .Q(n545) );
  INV6 U427 ( .A(n89), .Q(n524) );
  NAND23 U429 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND21 U430 ( .A(n556), .B(n51), .Q(n8) );
  NAND22 U433 ( .A(n111), .B(n554), .Q(n73) );
  INV1 U434 ( .A(n88), .Q(n562) );
  NAND21 U435 ( .A(n552), .B(n107), .Q(n14) );
  NAND24 U436 ( .A(B[24]), .B(A[24]), .Q(n107) );
  INV4 U437 ( .A(n97), .Q(n553) );
  AOI212 U439 ( .A(n523), .B(n97), .C(n98), .Q(n92) );
  NOR24 U440 ( .A(n46), .B(n6), .Q(n44) );
  NAND26 U441 ( .A(n524), .B(n525), .Q(n526) );
  NAND28 U442 ( .A(n436), .B(n437), .Q(SUM[30]) );
  NAND26 U443 ( .A(n532), .B(n555), .Q(n437) );
  AOI212 U444 ( .A(n523), .B(n554), .C(n551), .Q(n74) );
  NAND23 U445 ( .A(n517), .B(n518), .Q(n519) );
  NAND28 U446 ( .A(n519), .B(n100), .Q(n98) );
  CLKIN3 U448 ( .A(n99), .Q(n517) );
  INV6 U449 ( .A(n107), .Q(n518) );
  NAND22 U450 ( .A(B[11]), .B(A[11]), .Q(n224) );
  INV0 U452 ( .A(n513), .Q(n548) );
  NAND20 U453 ( .A(B[19]), .B(A[19]), .Q(n156) );
  OAI210 U454 ( .A(n126), .B(n543), .C(n127), .Q(n123) );
  INV0 U455 ( .A(n213), .Q(n572) );
  AOI210 U456 ( .A(n573), .B(n511), .C(n204), .Q(n198) );
  NAND21 U457 ( .A(n571), .B(n515), .Q(n26) );
  CLKIN6 U458 ( .A(n52), .Q(n532) );
  NAND21 U460 ( .A(n525), .B(n80), .Q(n11) );
  NAND22 U461 ( .A(B[27]), .B(A[27]), .Q(n80) );
  OAI211 U462 ( .A(n219), .B(n583), .C(n509), .Q(n214) );
  NAND22 U464 ( .A(n111), .B(n66), .Q(n64) );
  NOR22 U465 ( .A(n514), .B(n6), .Q(n66) );
  NOR24 U466 ( .A(n79), .B(n88), .Q(n77) );
  NAND22 U467 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NOR24 U468 ( .A(n61), .B(n70), .Q(n59) );
  AOI212 U471 ( .A(n523), .B(n84), .C(n85), .Q(n83) );
  NOR24 U472 ( .A(n99), .B(n106), .Q(n97) );
  NOR22 U473 ( .A(n260), .B(n265), .Q(n258) );
  BUF2 U474 ( .A(n117), .Q(n521) );
  INV2 U475 ( .A(n427), .Q(n551) );
  NAND22 U476 ( .A(n559), .B(n62), .Q(n9) );
  NAND22 U477 ( .A(A[29]), .B(B[29]), .Q(n62) );
  AOI210 U479 ( .A(n529), .B(n135), .C(n136), .Q(n130) );
  INV2 U480 ( .A(n152), .Q(n529) );
  INV1 U481 ( .A(n144), .Q(n549) );
  NAND24 U483 ( .A(n443), .B(n444), .Q(SUM[31]) );
  NAND24 U484 ( .A(n563), .B(n531), .Q(n444) );
  AOI212 U486 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  CLKIN1 U487 ( .A(n203), .Q(n569) );
  NOR24 U488 ( .A(n205), .B(n212), .Q(n203) );
  BUF15 U489 ( .A(n112), .Q(n523) );
  XNR22 U490 ( .A(n23), .B(n187), .Q(SUM[15]) );
  AOI212 U491 ( .A(n523), .B(n66), .C(n67), .Q(n65) );
  NOR24 U492 ( .A(n520), .B(n144), .Q(n135) );
  NAND22 U494 ( .A(n111), .B(n97), .Q(n91) );
  AOI212 U495 ( .A(n523), .B(n55), .C(n56), .Q(n54) );
  NAND22 U496 ( .A(A[9]), .B(B[9]), .Q(n242) );
  OAI211 U497 ( .A(n244), .B(n583), .C(n245), .Q(n243) );
  AOI210 U498 ( .A(n573), .B(n190), .C(n191), .Q(n189) );
  NOR21 U499 ( .A(n194), .B(n569), .Q(n190) );
  NAND23 U500 ( .A(A[16]), .B(B[16]), .Q(n177) );
  OAI212 U501 ( .A(n151), .B(n527), .C(n522), .Q(n146) );
  OAI212 U502 ( .A(n176), .B(n527), .C(n177), .Q(n175) );
  XNR22 U503 ( .A(n19), .B(n157), .Q(SUM[19]) );
  XNR22 U505 ( .A(n20), .B(n164), .Q(SUM[18]) );
  AOI210 U506 ( .A(n418), .B(n540), .C(n539), .Q(n159) );
  NAND20 U508 ( .A(n540), .B(n163), .Q(n20) );
  INV1 U509 ( .A(n162), .Q(n540) );
  XNR22 U510 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U512 ( .A(n15), .B(n119), .Q(SUM[23]) );
  OAI212 U514 ( .A(n64), .B(n527), .C(n65), .Q(n63) );
  NOR22 U515 ( .A(B[16]), .B(A[16]), .Q(n176) );
  XNR22 U516 ( .A(n17), .B(n139), .Q(SUM[21]) );
  OAI212 U517 ( .A(n152), .B(n113), .C(n114), .Q(n112) );
  OAI210 U518 ( .A(n173), .B(n177), .C(n174), .Q(n418) );
  NAND21 U519 ( .A(n549), .B(n513), .Q(n18) );
  XNR22 U521 ( .A(n18), .B(n146), .Q(SUM[20]) );
  INV2 U522 ( .A(n220), .Q(n573) );
  INV0 U523 ( .A(n512), .Q(n580) );
  XNR22 U524 ( .A(n21), .B(n175), .Q(SUM[17]) );
  XOR21 U525 ( .A(n32), .B(n257), .Q(SUM[6]) );
  OAI210 U526 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  XNR22 U527 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U528 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U529 ( .A(n12), .B(n90), .Q(SUM[26]) );
  XNR22 U530 ( .A(n11), .B(n81), .Q(SUM[27]) );
  CLKIN3 U532 ( .A(n6), .Q(n554) );
  NAND22 U533 ( .A(n111), .B(n55), .Q(n53) );
  NAND21 U534 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NOR22 U536 ( .A(n560), .B(n6), .Q(n55) );
  NAND22 U537 ( .A(n535), .B(n549), .Q(n140) );
  NAND28 U538 ( .A(n77), .B(n97), .Q(n6) );
  OAI211 U540 ( .A(n88), .B(n550), .C(n89), .Q(n85) );
  NAND22 U541 ( .A(B[21]), .B(A[21]), .Q(n138) );
  CLKIN2 U542 ( .A(n60), .Q(n558) );
  NAND21 U543 ( .A(n535), .B(n135), .Q(n129) );
  INV1 U544 ( .A(n219), .Q(n575) );
  INV1 U545 ( .A(n523), .Q(n530) );
  CLKIN0 U546 ( .A(n61), .Q(n559) );
  AOI212 U547 ( .A(n60), .B(n556), .C(n557), .Q(n47) );
  INV2 U548 ( .A(B[17]), .Q(n596) );
  INV0 U549 ( .A(n274), .Q(n590) );
  NAND20 U550 ( .A(n588), .B(n272), .Q(n35) );
  CLKIN6 U551 ( .A(n41), .Q(n531) );
  AOI212 U552 ( .A(n98), .B(n77), .C(n78), .Q(n427) );
  NAND20 U553 ( .A(n171), .B(n540), .Q(n158) );
  NAND20 U554 ( .A(n586), .B(n266), .Q(n34) );
  NAND20 U555 ( .A(n533), .B(n177), .Q(n22) );
  INV0 U556 ( .A(n176), .Q(n533) );
  NAND20 U557 ( .A(n584), .B(n256), .Q(n32) );
  NAND20 U558 ( .A(n590), .B(n275), .Q(n36) );
  NOR24 U559 ( .A(n252), .B(n255), .Q(n250) );
  AOI210 U560 ( .A(n573), .B(n571), .C(n572), .Q(n209) );
  INV0 U561 ( .A(n271), .Q(n588) );
  NAND20 U562 ( .A(n567), .B(n195), .Q(n24) );
  NOR24 U563 ( .A(n223), .B(n230), .Q(n221) );
  INV0 U564 ( .A(n266), .Q(n587) );
  NOR21 U565 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV2 U566 ( .A(A[17]), .Q(n537) );
  NOR22 U567 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND21 U568 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND21 U569 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND20 U570 ( .A(n592), .B(n279), .Q(n37) );
  INV0 U571 ( .A(n278), .Q(n592) );
  NAND21 U572 ( .A(A[31]), .B(B[31]), .Q(n40) );
  CLKIN3 U573 ( .A(n39), .Q(n564) );
  NAND22 U574 ( .A(n52), .B(n8), .Q(n436) );
  INV3 U575 ( .A(n8), .Q(n555) );
  NAND22 U576 ( .A(n575), .B(n511), .Q(n197) );
  NAND22 U577 ( .A(n575), .B(n190), .Q(n188) );
  NAND22 U578 ( .A(n575), .B(n571), .Q(n208) );
  NAND22 U579 ( .A(n122), .B(n535), .Q(n120) );
  INV3 U580 ( .A(n51), .Q(n557) );
  XOR20 U581 ( .A(n30), .B(n583), .Q(SUM[8]) );
  INV3 U582 ( .A(n244), .Q(n578) );
  INV3 U583 ( .A(n255), .Q(n584) );
  XOR21 U584 ( .A(n36), .B(n591), .Q(SUM[2]) );
  XNR21 U585 ( .A(n31), .B(n254), .Q(SUM[7]) );
  INV0 U586 ( .A(n252), .Q(n582) );
  XNR21 U587 ( .A(n35), .B(n273), .Q(SUM[3]) );
  INV0 U588 ( .A(n194), .Q(n567) );
  XNR21 U589 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND22 U590 ( .A(n574), .B(n224), .Q(n27) );
  INV0 U591 ( .A(n223), .Q(n574) );
  NAND20 U592 ( .A(n568), .B(n206), .Q(n25) );
  NAND22 U593 ( .A(n566), .B(n186), .Q(n23) );
  INV0 U594 ( .A(n185), .Q(n566) );
  XNR21 U595 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U596 ( .A(n576), .B(n231), .Q(n28) );
  XNR20 U597 ( .A(n34), .B(n589), .Q(SUM[4]) );
  NAND20 U598 ( .A(n174), .B(n538), .Q(n21) );
  INV0 U599 ( .A(n173), .Q(n538) );
  NAND22 U600 ( .A(n547), .B(n118), .Q(n15) );
  INV0 U601 ( .A(n521), .Q(n547) );
  NAND22 U602 ( .A(n542), .B(n156), .Q(n19) );
  INV0 U603 ( .A(n516), .Q(n542) );
  NAND22 U604 ( .A(n546), .B(n127), .Q(n16) );
  INV0 U605 ( .A(n126), .Q(n546) );
  NOR21 U606 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U607 ( .A(n258), .B(n250), .Q(n248) );
  NAND22 U608 ( .A(n581), .B(n242), .Q(n29) );
  INV0 U609 ( .A(n241), .Q(n581) );
  INV0 U610 ( .A(n99), .Q(n565) );
  INV0 U611 ( .A(n171), .Q(n534) );
  NAND22 U612 ( .A(n544), .B(n138), .Q(n17) );
  INV0 U613 ( .A(n520), .Q(n544) );
  XOR21 U614 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND22 U615 ( .A(n585), .B(n261), .Q(n33) );
  AOI210 U616 ( .A(n589), .B(n586), .C(n587), .Q(n262) );
  INV0 U617 ( .A(n260), .Q(n585) );
  NOR21 U618 ( .A(n126), .B(n545), .Q(n122) );
  AOI211 U619 ( .A(n529), .B(n122), .C(n123), .Q(n121) );
  AOI210 U620 ( .A(n512), .B(n576), .C(n577), .Q(n227) );
  INV0 U621 ( .A(n231), .Q(n577) );
  CLKIN1 U622 ( .A(n212), .Q(n571) );
  CLKIN0 U623 ( .A(n277), .Q(n591) );
  INV3 U624 ( .A(n230), .Q(n576) );
  CLKIN3 U625 ( .A(n106), .Q(n552) );
  INV3 U626 ( .A(n265), .Q(n586) );
  NOR21 U627 ( .A(n88), .B(n553), .Q(n84) );
  NAND22 U628 ( .A(n41), .B(n7), .Q(n443) );
  INV3 U629 ( .A(n7), .Q(n563) );
  XOR21 U630 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U631 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U632 ( .A(B[30]), .B(A[30]), .Q(n51) );
  NAND22 U633 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND22 U634 ( .A(B[6]), .B(A[6]), .Q(n256) );
  NAND22 U635 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U636 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND22 U637 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND22 U638 ( .A(n564), .B(n40), .Q(n7) );
  NOR21 U639 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U640 ( .A(A[0]), .B(B[0]), .Q(n281) );
  INV3 U641 ( .A(n38), .Q(SUM[0]) );
  NAND22 U642 ( .A(n594), .B(n281), .Q(n38) );
  INV3 U643 ( .A(n280), .Q(n594) );
  NOR21 U644 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U645 ( .A(n239), .B(n576), .Q(n226) );
  INV2 U646 ( .A(n239), .Q(n579) );
  OAI212 U647 ( .A(n5), .B(n560), .C(n558), .Q(n56) );
  NAND20 U648 ( .A(n562), .B(n89), .Q(n12) );
  CLKIN0 U649 ( .A(n514), .Q(n561) );
  NAND22 U650 ( .A(n561), .B(n71), .Q(n10) );
  NAND22 U651 ( .A(n565), .B(n100), .Q(n13) );
  CLKIN6 U652 ( .A(n79), .Q(n525) );
  NAND22 U653 ( .A(n111), .B(n552), .Q(n102) );
  NAND22 U654 ( .A(n111), .B(n84), .Q(n82) );
  INV2 U655 ( .A(n111), .Q(n536) );
  CLKIN0 U656 ( .A(n205), .Q(n568) );
  NAND20 U657 ( .A(B[17]), .B(A[17]), .Q(n174) );
  AOI212 U658 ( .A(n523), .B(n44), .C(n45), .Q(n43) );
endmodule


module adder_0 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1, n3, n4;

  adder_0_DW01_add_1 add_16 ( .A({A[31:22], n4, A[20:0]}), .B(B), .CI(n1), 
        .SUM(O) );
  CLKIN6 U1 ( .A(A[21]), .Q(n3) );
  INV12 U2 ( .A(n3), .Q(n4) );
  LOGIC0 U3 ( .Q(n1) );
endmodule


module reg_15 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n3, n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31,
         n34, n49, n51, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n108, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398;

  DF3 Dout_reg_14_ ( .D(n73), .C(Clk), .Q(Dout[14]), .QN(n3) );
  DF3 Dout_reg_13_ ( .D(n88), .C(Clk), .Q(Dout[13]), .QN(n78) );
  DF3 Dout_reg_12_ ( .D(n89), .C(Clk), .Q(Dout[12]), .QN(n74) );
  DF3 Dout_reg_11_ ( .D(n90), .C(Clk), .Q(Dout[11]), .QN(n76) );
  DF3 Dout_reg_10_ ( .D(n91), .C(Clk), .Q(Dout[10]), .QN(n75) );
  DF3 Dout_reg_9_ ( .D(n92), .C(Clk), .Q(Dout[9]), .QN(n77) );
  DF3 Dout_reg_8_ ( .D(n93), .C(Clk), .Q(Dout[8]), .QN(n79) );
  DF3 Dout_reg_7_ ( .D(n94), .C(Clk), .Q(Dout[7]), .QN(n82) );
  DF3 Dout_reg_6_ ( .D(n95), .C(Clk), .Q(Dout[6]), .QN(n81) );
  DF3 Dout_reg_5_ ( .D(n96), .C(Clk), .Q(Dout[5]), .QN(n80) );
  DF3 Dout_reg_4_ ( .D(n97), .C(Clk), .Q(Dout[4]), .QN(n84) );
  DF3 Dout_reg_3_ ( .D(n98), .C(Clk), .Q(Dout[3]), .QN(n85) );
  DF3 Dout_reg_2_ ( .D(n99), .C(Clk), .Q(Dout[2]), .QN(n83) );
  DF3 Dout_reg_1_ ( .D(n100), .C(Clk), .Q(Dout[1]), .QN(n87) );
  DF3 Dout_reg_0_ ( .D(n101), .C(Clk), .Q(Dout[0]), .QN(n86) );
  DF3 Dout_reg_15_ ( .D(n72), .C(Clk), .Q(Dout[15]), .QN(n5) );
  DF3 Dout_reg_16_ ( .D(n71), .C(Clk), .Q(Dout[16]), .QN(n7) );
  DF3 Dout_reg_17_ ( .D(n70), .C(Clk), .Q(Dout[17]), .QN(n9) );
  DF3 Dout_reg_18_ ( .D(n69), .C(Clk), .Q(Dout[18]), .QN(n11) );
  DF3 Dout_reg_24_ ( .D(n63), .C(Clk), .Q(Dout[24]), .QN(n23) );
  DF3 Dout_reg_22_ ( .D(n65), .C(Clk), .Q(Dout[22]), .QN(n19) );
  DF3 Dout_reg_19_ ( .D(n68), .C(Clk), .Q(Dout[19]), .QN(n13) );
  DF3 Dout_reg_20_ ( .D(n67), .C(Clk), .Q(Dout[20]), .QN(n15) );
  DF3 Dout_reg_21_ ( .D(n66), .C(Clk), .Q(Dout[21]), .QN(n17) );
  OAI222 U3 ( .A(n83), .B(n361), .C(n363), .D(n395), .Q(n99) );
  OAI222 U4 ( .A(n85), .B(n360), .C(n362), .D(n394), .Q(n98) );
  OAI222 U5 ( .A(n84), .B(n396), .C(n108), .D(n389), .Q(n97) );
  OAI222 U6 ( .A(n80), .B(n361), .C(n363), .D(n388), .Q(n96) );
  OAI222 U7 ( .A(n81), .B(n360), .C(n362), .D(n391), .Q(n95) );
  OAI222 U8 ( .A(n82), .B(n396), .C(n108), .D(n390), .Q(n94) );
  OAI222 U9 ( .A(n79), .B(n361), .C(n363), .D(n393), .Q(n93) );
  OAI222 U10 ( .A(n77), .B(n360), .C(n362), .D(n392), .Q(n92) );
  OAI222 U11 ( .A(n75), .B(n396), .C(n108), .D(n387), .Q(n91) );
  OAI222 U12 ( .A(n76), .B(n361), .C(n363), .D(n380), .Q(n90) );
  OAI222 U13 ( .A(n74), .B(n360), .C(n362), .D(n386), .Q(n89) );
  OAI222 U14 ( .A(n78), .B(n396), .C(n108), .D(n381), .Q(n88) );
  OAI222 U15 ( .A(n3), .B(n361), .C(n363), .D(n382), .Q(n73) );
  OAI222 U16 ( .A(n5), .B(n360), .C(n362), .D(n383), .Q(n72) );
  OAI222 U17 ( .A(n7), .B(n396), .C(n108), .D(n384), .Q(n71) );
  OAI222 U18 ( .A(n9), .B(n361), .C(n385), .D(n363), .Q(n70) );
  OAI222 U19 ( .A(n11), .B(n360), .C(n379), .D(n362), .Q(n69) );
  OAI222 U20 ( .A(n13), .B(n396), .C(n378), .D(n108), .Q(n68) );
  OAI222 U21 ( .A(n15), .B(n361), .C(n377), .D(n363), .Q(n67) );
  OAI222 U22 ( .A(n17), .B(n360), .C(n376), .D(n362), .Q(n66) );
  OAI222 U23 ( .A(n19), .B(n396), .C(n375), .D(n108), .Q(n65) );
  OAI222 U24 ( .A(n21), .B(n361), .C(n374), .D(n363), .Q(n64) );
  OAI222 U25 ( .A(n23), .B(n360), .C(n373), .D(n362), .Q(n63) );
  OAI222 U26 ( .A(n25), .B(n396), .C(n372), .D(n108), .Q(n62) );
  OAI222 U27 ( .A(n27), .B(n361), .C(n371), .D(n363), .Q(n61) );
  OAI222 U28 ( .A(n29), .B(n360), .C(n370), .D(n362), .Q(n60) );
  OAI222 U29 ( .A(n31), .B(n396), .C(n369), .D(n108), .Q(n59) );
  OAI222 U31 ( .A(n49), .B(n361), .C(n368), .D(n363), .Q(n57) );
  OAI222 U32 ( .A(n51), .B(n360), .C(n367), .D(n362), .Q(n56) );
  OAI222 U33 ( .A(n86), .B(n396), .C(n108), .D(n398), .Q(n101) );
  OAI222 U34 ( .A(n87), .B(n361), .C(n363), .D(n397), .Q(n100) );
  DF1 Dout_reg_28_ ( .D(n59), .C(Clk), .Q(Dout[28]), .QN(n31) );
  DF1 Dout_reg_27_ ( .D(n60), .C(Clk), .Q(Dout[27]), .QN(n29) );
  DF1 Dout_reg_31_ ( .D(n56), .C(Clk), .Q(Dout[31]), .QN(n51) );
  DF1 Dout_reg_30_ ( .D(n57), .C(Clk), .Q(Dout[30]), .QN(n49) );
  DF1 Dout_reg_25_ ( .D(n62), .C(Clk), .Q(Dout[25]), .QN(n25) );
  DF1 Dout_reg_29_ ( .D(n58), .C(Clk), .Q(Dout[29]), .QN(n34) );
  DF3 Dout_reg_26_ ( .D(n61), .C(Clk), .Q(Dout[26]), .QN(n27) );
  DF1 Dout_reg_23_ ( .D(n64), .C(Clk), .Q(Dout[23]), .QN(n21) );
  INV4 U30 ( .A(Din[31]), .Q(n367) );
  INV4 U35 ( .A(Din[26]), .Q(n371) );
  INV4 U36 ( .A(Din[25]), .Q(n372) );
  INV2 U37 ( .A(Din[16]), .Q(n384) );
  INV2 U38 ( .A(Din[12]), .Q(n386) );
  INV4 U39 ( .A(Din[20]), .Q(n377) );
  INV4 U40 ( .A(Din[17]), .Q(n385) );
  INV4 U41 ( .A(Din[22]), .Q(n375) );
  INV3 U42 ( .A(Din[15]), .Q(n383) );
  INV4 U43 ( .A(Din[24]), .Q(n373) );
  INV4 U44 ( .A(Din[21]), .Q(n376) );
  INV4 U45 ( .A(Din[23]), .Q(n374) );
  INV4 U46 ( .A(Din[18]), .Q(n379) );
  INV4 U47 ( .A(Din[19]), .Q(n378) );
  INV4 U48 ( .A(Din[28]), .Q(n369) );
  INV4 U49 ( .A(Din[27]), .Q(n370) );
  INV4 U50 ( .A(Din[30]), .Q(n368) );
  INV3 U51 ( .A(Din[29]), .Q(n366) );
  INV2 U52 ( .A(Din[14]), .Q(n382) );
  INV2 U53 ( .A(Din[13]), .Q(n381) );
  INV2 U54 ( .A(Din[11]), .Q(n380) );
  INV2 U55 ( .A(Din[9]), .Q(n392) );
  CLKIN2 U56 ( .A(Din[8]), .Q(n393) );
  INV2 U57 ( .A(Din[10]), .Q(n387) );
  INV3 U58 ( .A(Reset), .Q(n364) );
  NAND22 U59 ( .A(n364), .B(n365), .Q(n360) );
  NAND22 U60 ( .A(n364), .B(n365), .Q(n361) );
  NAND22 U61 ( .A(n364), .B(n365), .Q(n396) );
  INV3 U62 ( .A(Din[7]), .Q(n390) );
  INV3 U63 ( .A(Din[6]), .Q(n391) );
  INV3 U64 ( .A(Din[2]), .Q(n395) );
  INV3 U65 ( .A(Din[3]), .Q(n394) );
  INV3 U66 ( .A(Din[5]), .Q(n388) );
  INV3 U67 ( .A(Din[4]), .Q(n389) );
  NAND22 U68 ( .A(Load), .B(n364), .Q(n362) );
  NAND22 U69 ( .A(Load), .B(n364), .Q(n363) );
  NAND22 U70 ( .A(Load), .B(n364), .Q(n108) );
  INV3 U71 ( .A(Din[1]), .Q(n397) );
  INV3 U72 ( .A(Din[0]), .Q(n398) );
  INV1 U73 ( .A(Load), .Q(n365) );
  OAI222 U74 ( .A(n34), .B(n360), .C(n366), .D(n362), .Q(n58) );
endmodule


module reg_14 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30,
         n32, n35, n47, n49, n51, n53, n55, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n58, n59, n60, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n102, n103, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393;

  DF3 Dout_reg_16_ ( .D(n76), .C(Clk), .Q(Dout[16]), .QN(n14) );
  DF3 Dout_reg_15_ ( .D(n77), .C(Clk), .Q(Dout[15]), .QN(n12) );
  DF3 Dout_reg_14_ ( .D(n78), .C(Clk), .Q(Dout[14]), .QN(n10) );
  DF3 Dout_reg_13_ ( .D(n79), .C(Clk), .Q(Dout[13]), .QN(n8) );
  DF3 Dout_reg_12_ ( .D(n80), .C(Clk), .Q(Dout[12]), .QN(n6) );
  DF3 Dout_reg_11_ ( .D(n81), .C(Clk), .Q(Dout[11]), .QN(n4) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n82) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n59) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n58) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n86) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n83) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n85) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n84) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n87) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n88) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n89) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n60) );
  OAI222 U3 ( .A(n88), .B(n358), .C(n360), .D(n392), .Q(n99) );
  OAI222 U4 ( .A(n87), .B(n358), .C(n359), .D(n391), .Q(n98) );
  OAI222 U5 ( .A(n84), .B(n358), .C(n102), .D(n390), .Q(n97) );
  OAI222 U6 ( .A(n85), .B(n358), .C(n360), .D(n389), .Q(n96) );
  OAI222 U7 ( .A(n83), .B(n358), .C(n359), .D(n388), .Q(n95) );
  OAI222 U8 ( .A(n86), .B(n358), .C(n102), .D(n387), .Q(n94) );
  OAI222 U9 ( .A(n58), .B(n358), .C(n360), .D(n386), .Q(n93) );
  OAI222 U10 ( .A(n59), .B(n358), .C(n359), .D(n385), .Q(n92) );
  OAI222 U11 ( .A(n60), .B(n358), .C(n102), .D(n384), .Q(n91) );
  OAI222 U12 ( .A(n82), .B(n358), .C(n360), .D(n383), .Q(n90) );
  OAI222 U13 ( .A(n4), .B(n358), .C(n359), .D(n382), .Q(n81) );
  OAI222 U14 ( .A(n6), .B(n358), .C(n102), .D(n381), .Q(n80) );
  OAI222 U15 ( .A(n8), .B(n358), .C(n360), .D(n380), .Q(n79) );
  OAI222 U16 ( .A(n10), .B(n358), .C(n359), .D(n379), .Q(n78) );
  OAI222 U17 ( .A(n12), .B(n358), .C(n102), .D(n378), .Q(n77) );
  OAI222 U18 ( .A(n14), .B(n358), .C(n360), .D(n374), .Q(n76) );
  OAI222 U19 ( .A(n16), .B(n358), .C(n359), .D(n377), .Q(n75) );
  OAI222 U20 ( .A(n18), .B(n358), .C(n102), .D(n375), .Q(n74) );
  OAI222 U21 ( .A(n20), .B(n358), .C(n360), .D(n376), .Q(n73) );
  OAI222 U22 ( .A(n22), .B(n358), .C(n359), .D(n365), .Q(n72) );
  OAI222 U23 ( .A(n24), .B(n358), .C(n363), .D(n102), .Q(n71) );
  OAI222 U24 ( .A(n26), .B(n358), .C(n360), .D(n362), .Q(n70) );
  OAI222 U25 ( .A(n28), .B(n358), .C(n359), .D(n364), .Q(n69) );
  OAI222 U26 ( .A(n30), .B(n358), .C(n102), .D(n372), .Q(n68) );
  OAI222 U27 ( .A(n32), .B(n358), .C(n360), .D(n368), .Q(n67) );
  OAI222 U28 ( .A(n35), .B(n358), .C(n359), .D(n373), .Q(n66) );
  OAI222 U29 ( .A(n47), .B(n358), .C(n102), .D(n367), .Q(n65) );
  OAI222 U30 ( .A(n49), .B(n358), .C(n369), .D(n360), .Q(n64) );
  OAI222 U31 ( .A(n51), .B(n358), .C(n370), .D(n359), .Q(n63) );
  OAI222 U32 ( .A(n53), .B(n358), .C(n102), .D(n366), .Q(n62) );
  OAI222 U33 ( .A(n55), .B(n358), .C(n360), .D(n371), .Q(n61) );
  OAI222 U34 ( .A(n89), .B(n358), .C(n359), .D(n393), .Q(n100) );
  DF1 Dout_reg_30_ ( .D(n62), .C(Clk), .Q(Dout[30]), .QN(n53) );
  DF1 Dout_reg_31_ ( .D(n61), .C(Clk), .Q(Dout[31]), .QN(n55) );
  DF1 Dout_reg_28_ ( .D(n64), .C(Clk), .Q(Dout[28]), .QN(n49) );
  DF1 Dout_reg_22_ ( .D(n70), .C(Clk), .Q(Dout[22]), .QN(n26) );
  DF1 Dout_reg_21_ ( .D(n71), .C(Clk), .Q(Dout[21]), .QN(n24) );
  DF1 Dout_reg_20_ ( .D(n72), .C(Clk), .Q(Dout[20]), .QN(n22) );
  DF1 Dout_reg_18_ ( .D(n74), .C(Clk), .Q(Dout[18]), .QN(n18) );
  DF1 Dout_reg_26_ ( .D(n66), .C(Clk), .Q(Dout[26]), .QN(n35) );
  DF1 Dout_reg_27_ ( .D(n65), .C(Clk), .Q(Dout[27]), .QN(n47) );
  DF1 Dout_reg_17_ ( .D(n75), .C(Clk), .Q(Dout[17]), .QN(n16) );
  DF3 Dout_reg_23_ ( .D(n69), .C(Clk), .Q(Dout[23]), .QN(n28) );
  DF3 Dout_reg_24_ ( .D(n68), .C(Clk), .Q(Dout[24]), .QN(n30) );
  DF3 Dout_reg_19_ ( .D(n73), .C(Clk), .Q(Dout[19]), .QN(n20) );
  DF1 Dout_reg_29_ ( .D(n63), .C(Clk), .Q(Dout[29]), .QN(n51) );
  DF1 Dout_reg_25_ ( .D(n67), .C(Clk), .Q(Dout[25]), .QN(n32) );
  INV3 U35 ( .A(Din[29]), .Q(n370) );
  CLKIN6 U36 ( .A(Din[26]), .Q(n373) );
  INV3 U37 ( .A(Din[17]), .Q(n377) );
  INV3 U38 ( .A(Din[20]), .Q(n365) );
  INV3 U39 ( .A(Din[24]), .Q(n372) );
  INV3 U40 ( .A(Din[31]), .Q(n371) );
  INV3 U41 ( .A(Din[28]), .Q(n369) );
  INV3 U42 ( .A(Din[30]), .Q(n366) );
  CLKIN3 U43 ( .A(Din[7]), .Q(n386) );
  INV2 U44 ( .A(Din[15]), .Q(n378) );
  INV2 U45 ( .A(Din[14]), .Q(n379) );
  INV2 U46 ( .A(Din[13]), .Q(n380) );
  CLKIN3 U47 ( .A(Din[8]), .Q(n385) );
  INV2 U48 ( .A(Din[6]), .Q(n387) );
  INV2 U49 ( .A(Din[25]), .Q(n368) );
  INV2 U50 ( .A(Din[23]), .Q(n364) );
  INV2 U51 ( .A(Din[22]), .Q(n362) );
  INV2 U52 ( .A(Din[27]), .Q(n367) );
  INV2 U53 ( .A(Din[21]), .Q(n363) );
  INV2 U54 ( .A(Din[19]), .Q(n376) );
  INV2 U55 ( .A(Din[16]), .Q(n374) );
  INV2 U56 ( .A(Din[11]), .Q(n382) );
  INV2 U57 ( .A(Din[10]), .Q(n383) );
  INV2 U58 ( .A(Din[18]), .Q(n375) );
  INV2 U59 ( .A(Din[12]), .Q(n381) );
  INV2 U60 ( .A(Din[9]), .Q(n384) );
  NAND22 U61 ( .A(n361), .B(n358), .Q(n359) );
  NAND22 U62 ( .A(n361), .B(n358), .Q(n360) );
  NAND22 U63 ( .A(n361), .B(n358), .Q(n102) );
  INV3 U64 ( .A(Reset), .Q(n361) );
  INV3 U65 ( .A(n103), .Q(n358) );
  INV3 U66 ( .A(Din[4]), .Q(n389) );
  INV3 U67 ( .A(Din[5]), .Q(n388) );
  INV3 U68 ( .A(Din[1]), .Q(n392) );
  INV3 U69 ( .A(Din[3]), .Q(n390) );
  INV3 U70 ( .A(Din[2]), .Q(n391) );
  INV3 U71 ( .A(Din[0]), .Q(n393) );
  NOR20 U72 ( .A(Load), .B(Reset), .Q(n103) );
endmodule


module adder_45_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n416, n417,
         n551, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816;

  OAI212 U15 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U43 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI212 U51 ( .A(n73), .B(n753), .C(n74), .Q(n72) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n753), .C(n121), .Q(n119) );
  OAI212 U127 ( .A(n129), .B(n753), .C(n130), .Q(n128) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n753), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U159 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U165 ( .A(n158), .B(n753), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n758), .B(n753), .C(n754), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n777), .C(n227), .Q(n225) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  AOI212 U371 ( .A(n277), .B(n269), .C(n270), .Q(n416) );
  OAI212 U375 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U376 ( .A(n248), .B(n268), .C(n249), .Q(n417) );
  OAI212 U354 ( .A(n775), .B(n777), .C(n773), .Q(n232) );
  OAI212 U358 ( .A(n760), .B(n753), .C(n756), .Q(n108) );
  OAI212 U433 ( .A(n208), .B(n777), .C(n209), .Q(n207) );
  OAI212 U360 ( .A(n188), .B(n777), .C(n189), .Q(n187) );
  OAI212 U427 ( .A(n248), .B(n416), .C(n249), .Q(n247) );
  OAI212 U442 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U351 ( .A(n194), .B(n765), .C(n195), .Q(n191) );
  OAI212 U423 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NOR24 U356 ( .A(B[3]), .B(A[3]), .Q(n271) );
  OAI212 U399 ( .A(n244), .B(n777), .C(n245), .Q(n243) );
  OAI212 U402 ( .A(n102), .B(n753), .C(n103), .Q(n101) );
  OAI212 U409 ( .A(n176), .B(n753), .C(n177), .Q(n175) );
  OAI212 U406 ( .A(n42), .B(n753), .C(n43), .Q(n41) );
  OAI212 U431 ( .A(n53), .B(n753), .C(n54), .Q(n52) );
  OAI212 U499 ( .A(n795), .B(n5), .C(n793), .Q(n56) );
  NOR24 U389 ( .A(B[9]), .B(A[9]), .Q(n241) );
  XNR22 U392 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U407 ( .A(n23), .B(n187), .Q(SUM[15]) );
  OAI212 U411 ( .A(n82), .B(n753), .C(n83), .Q(n81) );
  AOI212 U413 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  XNR22 U425 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR22 U426 ( .A(n15), .B(n119), .Q(SUM[23]) );
  XNR22 U428 ( .A(n29), .B(n243), .Q(SUM[9]) );
  XNR22 U429 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U432 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U438 ( .A(n12), .B(n90), .Q(SUM[26]) );
  XNR22 U439 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U441 ( .A(n27), .B(n225), .Q(SUM[11]) );
  XNR22 U447 ( .A(n20), .B(n164), .Q(SUM[18]) );
  XNR22 U450 ( .A(n19), .B(n157), .Q(SUM[19]) );
  XNR22 U451 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NOR24 U350 ( .A(n185), .B(n194), .Q(n183) );
  OAI212 U366 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U391 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U436 ( .A(n64), .B(n753), .C(n65), .Q(n63) );
  OAI212 U443 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NOR24 U449 ( .A(B[10]), .B(A[10]), .Q(n230) );
  OAI212 U465 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U466 ( .A(n88), .B(n800), .C(n89), .Q(n85) );
  XOR22 U561 ( .A(n33), .B(n752), .Q(SUM[5]) );
  XNR22 U565 ( .A(n24), .B(n196), .Q(SUM[14]) );
  XNR22 U579 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U584 ( .A(n10), .B(n72), .Q(SUM[28]) );
  INV2 U349 ( .A(n262), .Q(n751) );
  NAND22 U352 ( .A(n111), .B(n55), .Q(n53) );
  NAND22 U353 ( .A(n111), .B(n797), .Q(n102) );
  NOR23 U355 ( .A(n223), .B(n230), .Q(n221) );
  NOR23 U357 ( .A(B[11]), .B(A[11]), .Q(n223) );
  INV2 U359 ( .A(n220), .Q(n768) );
  BUF15 U361 ( .A(n178), .Q(n753) );
  NOR23 U362 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND28 U363 ( .A(n239), .B(n221), .Q(n219) );
  NOR22 U364 ( .A(n241), .B(n244), .Q(n239) );
  XOR22 U365 ( .A(n22), .B(n753), .Q(SUM[16]) );
  XNR22 U367 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND22 U368 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NOR23 U369 ( .A(n252), .B(n255), .Q(n250) );
  NOR23 U370 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR22 U372 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR22 U373 ( .A(n79), .B(n88), .Q(n77) );
  NOR22 U374 ( .A(n117), .B(n126), .Q(n115) );
  NOR21 U377 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR21 U378 ( .A(B[24]), .B(A[24]), .Q(n106) );
  XNR21 U379 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NOR22 U380 ( .A(B[7]), .B(A[7]), .Q(n252) );
  INV3 U381 ( .A(n416), .Q(n782) );
  AOI211 U382 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  INV6 U383 ( .A(n417), .Q(n777) );
  NOR23 U384 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NAND22 U385 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NOR22 U386 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR22 U387 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U388 ( .A(n88), .B(n798), .Q(n84) );
  AOI211 U390 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  AOI211 U393 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NOR21 U394 ( .A(n70), .B(n6), .Q(n66) );
  XNR21 U395 ( .A(n26), .B(n214), .Q(SUM[12]) );
  AOI211 U396 ( .A(n755), .B(n803), .C(n805), .Q(n141) );
  NOR22 U397 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND22 U398 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NOR23 U400 ( .A(n113), .B(n151), .Q(n111) );
  NAND22 U401 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NOR22 U403 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR22 U404 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR22 U405 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR22 U408 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR22 U410 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR23 U412 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR22 U414 ( .A(B[1]), .B(A[1]), .Q(n278) );
  XNR21 U415 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XNR21 U416 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NOR22 U417 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR21 U418 ( .A(n181), .B(n219), .Q(n179) );
  XOR21 U419 ( .A(n30), .B(n777), .Q(SUM[8]) );
  XOR21 U420 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND22 U421 ( .A(A[0]), .B(B[0]), .Q(n281) );
  INV3 U422 ( .A(n112), .Q(n756) );
  INV3 U424 ( .A(n751), .Q(n752) );
  AOI212 U430 ( .A(n112), .B(n97), .C(n98), .Q(n92) );
  NOR22 U434 ( .A(n155), .B(n162), .Q(n153) );
  OAI211 U435 ( .A(n91), .B(n753), .C(n92), .Q(n90) );
  INV1 U437 ( .A(n277), .Q(n785) );
  NOR23 U440 ( .A(n271), .B(n274), .Q(n269) );
  INV2 U444 ( .A(n151), .Q(n759) );
  AOI211 U445 ( .A(n768), .B(n203), .C(n204), .Q(n198) );
  NOR22 U446 ( .A(n99), .B(n106), .Q(n97) );
  NOR22 U448 ( .A(B[25]), .B(A[25]), .Q(n99) );
  AOI211 U452 ( .A(n755), .B(n122), .C(n123), .Q(n121) );
  NAND21 U453 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NOR22 U454 ( .A(n173), .B(n176), .Q(n171) );
  NOR22 U455 ( .A(B[17]), .B(A[17]), .Q(n173) );
  OAI211 U456 ( .A(n275), .B(n271), .C(n272), .Q(n551) );
  AOI212 U457 ( .A(n112), .B(n797), .C(n799), .Q(n103) );
  NAND21 U458 ( .A(n810), .B(n156), .Q(n19) );
  OAI211 U459 ( .A(n197), .B(n777), .C(n198), .Q(n196) );
  INV3 U460 ( .A(n219), .Q(n770) );
  AOI211 U461 ( .A(n84), .B(n112), .C(n85), .Q(n83) );
  INV1 U462 ( .A(n135), .Q(n804) );
  AOI211 U463 ( .A(n755), .B(n135), .C(n136), .Q(n130) );
  NAND23 U464 ( .A(n135), .B(n115), .Q(n113) );
  NAND22 U467 ( .A(n759), .B(n135), .Q(n129) );
  NOR23 U468 ( .A(n137), .B(n144), .Q(n135) );
  NOR21 U469 ( .A(n126), .B(n804), .Q(n122) );
  NAND24 U470 ( .A(A[8]), .B(B[8]), .Q(n245) );
  XNR22 U471 ( .A(n18), .B(n146), .Q(SUM[20]) );
  OAI211 U472 ( .A(n151), .B(n753), .C(n152), .Q(n146) );
  AOI212 U473 ( .A(n782), .B(n258), .C(n259), .Q(n257) );
  XOR20 U474 ( .A(n36), .B(n785), .Q(SUM[2]) );
  OAI211 U475 ( .A(n274), .B(n785), .C(n275), .Q(n273) );
  OAI211 U476 ( .A(n219), .B(n777), .C(n220), .Q(n214) );
  INV2 U477 ( .A(n152), .Q(n755) );
  NAND20 U478 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND21 U479 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NAND21 U480 ( .A(n797), .B(n107), .Q(n14) );
  INV2 U481 ( .A(n6), .Q(n792) );
  INV1 U482 ( .A(n111), .Q(n760) );
  NAND23 U483 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U484 ( .A(n791), .B(n89), .Q(n12) );
  INV0 U485 ( .A(n88), .Q(n791) );
  NAND20 U486 ( .A(n796), .B(n80), .Q(n11) );
  NAND21 U487 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND20 U488 ( .A(n770), .B(n203), .Q(n197) );
  NAND23 U489 ( .A(n258), .B(n250), .Q(n248) );
  INV0 U490 ( .A(n230), .Q(n771) );
  NAND20 U491 ( .A(n769), .B(n224), .Q(n27) );
  NAND20 U492 ( .A(n803), .B(n145), .Q(n18) );
  NAND21 U493 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NAND21 U494 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND22 U495 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NOR20 U496 ( .A(n795), .B(n6), .Q(n55) );
  NAND21 U497 ( .A(n770), .B(n190), .Q(n188) );
  CLKIN3 U498 ( .A(n59), .Q(n795) );
  INV0 U500 ( .A(n99), .Q(n811) );
  NAND20 U501 ( .A(n811), .B(n100), .Q(n13) );
  INV0 U502 ( .A(n79), .Q(n796) );
  NAND20 U503 ( .A(n783), .B(n272), .Q(n35) );
  XOR20 U504 ( .A(n281), .B(n37), .Q(SUM[1]) );
  XNR20 U505 ( .A(n34), .B(n782), .Q(SUM[4]) );
  NAND20 U506 ( .A(n780), .B(n266), .Q(n34) );
  NOR20 U507 ( .A(n194), .B(n764), .Q(n190) );
  NOR23 U508 ( .A(n205), .B(n212), .Q(n203) );
  INV0 U509 ( .A(n173), .Q(n809) );
  NAND20 U510 ( .A(n779), .B(n261), .Q(n33) );
  AOI210 U511 ( .A(n782), .B(n780), .C(n781), .Q(n262) );
  INV0 U512 ( .A(n126), .Q(n807) );
  INV0 U513 ( .A(n241), .Q(n789) );
  NAND20 U514 ( .A(n789), .B(n242), .Q(n29) );
  OAI211 U515 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND20 U516 ( .A(n762), .B(n195), .Q(n24) );
  INV1 U517 ( .A(n61), .Q(n815) );
  INV0 U518 ( .A(n117), .Q(n808) );
  CLKIN1 U519 ( .A(n106), .Q(n797) );
  NAND21 U520 ( .A(n59), .B(n813), .Q(n46) );
  OAI210 U521 ( .A(n126), .B(n806), .C(n127), .Q(n123) );
  INV0 U522 ( .A(n266), .Q(n781) );
  NOR22 U523 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR22 U524 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR22 U525 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NAND21 U526 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND21 U527 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NAND21 U528 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND21 U529 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND21 U530 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND21 U531 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND22 U532 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND22 U533 ( .A(n111), .B(n792), .Q(n73) );
  NAND20 U534 ( .A(n111), .B(n44), .Q(n42) );
  AOI210 U535 ( .A(n112), .B(n792), .C(n790), .Q(n74) );
  CLKIN1 U536 ( .A(n5), .Q(n790) );
  AOI210 U537 ( .A(n112), .B(n55), .C(n56), .Q(n54) );
  INV3 U538 ( .A(n60), .Q(n793) );
  NAND22 U539 ( .A(n97), .B(n77), .Q(n6) );
  NOR20 U540 ( .A(n46), .B(n6), .Q(n44) );
  NAND22 U541 ( .A(n171), .B(n153), .Q(n151) );
  NAND20 U542 ( .A(n111), .B(n84), .Q(n82) );
  NAND20 U543 ( .A(n111), .B(n66), .Q(n64) );
  NAND20 U544 ( .A(n111), .B(n97), .Q(n91) );
  NAND24 U545 ( .A(n203), .B(n183), .Q(n181) );
  NAND20 U546 ( .A(n239), .B(n771), .Q(n226) );
  INV0 U547 ( .A(n239), .Q(n775) );
  NAND22 U548 ( .A(n759), .B(n122), .Q(n120) );
  NAND22 U549 ( .A(n759), .B(n803), .Q(n140) );
  NAND22 U550 ( .A(n171), .B(n801), .Q(n158) );
  NAND22 U551 ( .A(n770), .B(n766), .Q(n208) );
  INV0 U552 ( .A(n172), .Q(n754) );
  NAND22 U553 ( .A(n815), .B(n62), .Q(n9) );
  INV3 U554 ( .A(n107), .Q(n799) );
  INV0 U555 ( .A(n98), .Q(n800) );
  AOI210 U556 ( .A(n112), .B(n66), .C(n67), .Q(n65) );
  NAND22 U557 ( .A(n778), .B(n256), .Q(n32) );
  INV0 U558 ( .A(n255), .Q(n778) );
  NAND22 U559 ( .A(n813), .B(n51), .Q(n8) );
  NAND22 U560 ( .A(n807), .B(n127), .Q(n16) );
  NAND22 U562 ( .A(n786), .B(n279), .Q(n37) );
  INV0 U563 ( .A(n278), .Q(n786) );
  NAND22 U564 ( .A(n757), .B(n177), .Q(n22) );
  INV3 U566 ( .A(n176), .Q(n757) );
  INV0 U567 ( .A(n260), .Q(n779) );
  NAND22 U568 ( .A(n774), .B(n245), .Q(n30) );
  INV0 U569 ( .A(n244), .Q(n774) );
  NAND22 U570 ( .A(n784), .B(n275), .Q(n36) );
  INV3 U571 ( .A(n274), .Q(n784) );
  INV3 U572 ( .A(n231), .Q(n772) );
  XNR21 U573 ( .A(n35), .B(n273), .Q(SUM[3]) );
  INV0 U574 ( .A(n271), .Q(n783) );
  NAND22 U575 ( .A(n761), .B(n186), .Q(n23) );
  INV0 U576 ( .A(n185), .Q(n761) );
  INV0 U577 ( .A(n194), .Q(n762) );
  NAND22 U578 ( .A(n809), .B(n174), .Q(n21) );
  NAND22 U580 ( .A(n766), .B(n213), .Q(n26) );
  INV3 U581 ( .A(n155), .Q(n810) );
  NAND22 U582 ( .A(n812), .B(n138), .Q(n17) );
  INV3 U583 ( .A(n137), .Q(n812) );
  NOR21 U585 ( .A(n61), .B(n70), .Q(n59) );
  NAND22 U586 ( .A(n794), .B(n71), .Q(n10) );
  INV3 U587 ( .A(n70), .Q(n794) );
  AOI210 U588 ( .A(n112), .B(n44), .C(n45), .Q(n43) );
  AOI211 U589 ( .A(n60), .B(n813), .C(n814), .Q(n47) );
  INV3 U590 ( .A(n51), .Q(n814) );
  NAND22 U591 ( .A(n776), .B(n253), .Q(n31) );
  INV0 U592 ( .A(n252), .Q(n776) );
  CLKIN0 U593 ( .A(n223), .Q(n769) );
  NAND22 U594 ( .A(n771), .B(n231), .Q(n28) );
  INV0 U595 ( .A(n240), .Q(n773) );
  NAND22 U596 ( .A(n808), .B(n118), .Q(n15) );
  NAND22 U597 ( .A(n801), .B(n163), .Q(n20) );
  INV0 U598 ( .A(n171), .Q(n758) );
  INV3 U599 ( .A(n97), .Q(n798) );
  NAND22 U600 ( .A(n763), .B(n206), .Q(n25) );
  INV0 U601 ( .A(n205), .Q(n763) );
  NOR22 U602 ( .A(n260), .B(n265), .Q(n258) );
  AOI210 U603 ( .A(n172), .B(n801), .C(n802), .Q(n159) );
  INV3 U604 ( .A(n163), .Q(n802) );
  INV0 U605 ( .A(n136), .Q(n806) );
  AOI211 U606 ( .A(n768), .B(n190), .C(n191), .Q(n189) );
  INV0 U607 ( .A(n204), .Q(n765) );
  INV3 U608 ( .A(n145), .Q(n805) );
  AOI211 U609 ( .A(n768), .B(n766), .C(n767), .Q(n209) );
  INV3 U610 ( .A(n213), .Q(n767) );
  INV3 U611 ( .A(n144), .Q(n803) );
  INV3 U612 ( .A(n162), .Q(n801) );
  CLKIN1 U613 ( .A(n212), .Q(n766) );
  INV1 U614 ( .A(n203), .Q(n764) );
  CLKIN0 U615 ( .A(n265), .Q(n780) );
  NOR22 U616 ( .A(B[28]), .B(A[28]), .Q(n70) );
  XNR21 U617 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U618 ( .A(n816), .B(n40), .Q(n7) );
  NAND22 U619 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR21 U620 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND22 U621 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND22 U622 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND22 U623 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND21 U624 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND21 U625 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND22 U626 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND22 U627 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND22 U628 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U629 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV3 U630 ( .A(n50), .Q(n813) );
  NOR21 U631 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U632 ( .A(n38), .Q(SUM[0]) );
  NAND20 U633 ( .A(n788), .B(n281), .Q(n38) );
  INV3 U634 ( .A(n280), .Q(n788) );
  NOR20 U635 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U636 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U637 ( .A(n39), .Q(n816) );
  NOR21 U638 ( .A(B[31]), .B(A[31]), .Q(n39) );
  AOI211 U639 ( .A(n277), .B(n269), .C(n551), .Q(n268) );
  AOI210 U640 ( .A(n240), .B(n771), .C(n772), .Q(n227) );
endmodule


module adder_45 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_45_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_44_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n50,
         n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n416, n417, n419,
         n420, n423, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n508, n509, n510;

  OAI212 U11 ( .A(n42), .B(n444), .C(n43), .Q(n41) );
  OAI212 U25 ( .A(n53), .B(n444), .C(n54), .Q(n52) );
  OAI212 U65 ( .A(n82), .B(n444), .C(n83), .Q(n81) );
  OAI212 U101 ( .A(n444), .B(n465), .C(n463), .Q(n108) );
  OAI212 U115 ( .A(n120), .B(n444), .C(n121), .Q(n119) );
  OAI212 U127 ( .A(n129), .B(n444), .C(n130), .Q(n128) );
  OAI212 U141 ( .A(n140), .B(n444), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U159 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U165 ( .A(n158), .B(n444), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n490), .B(n444), .C(n488), .Q(n164) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U219 ( .A(n197), .B(n495), .C(n198), .Q(n196) );
  OAI212 U227 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  OAI212 U233 ( .A(n208), .B(n495), .C(n209), .Q(n207) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U257 ( .A(n226), .B(n495), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n499), .B(n495), .C(n500), .Q(n232) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n508), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U491 ( .A(n73), .B(n444), .C(n74), .Q(n72) );
  OAI212 U494 ( .A(n444), .B(n102), .C(n103), .Q(n101) );
  OAI212 U403 ( .A(n88), .B(n456), .C(n89), .Q(n85) );
  NAND22 U349 ( .A(n100), .B(n457), .Q(n13) );
  INV1 U350 ( .A(n203), .Q(n482) );
  NAND21 U351 ( .A(n111), .B(n97), .Q(n91) );
  INV2 U352 ( .A(n499), .Q(n428) );
  INV3 U353 ( .A(n239), .Q(n499) );
  OAI211 U354 ( .A(n252), .B(n256), .C(n253), .Q(n251) );
  NAND26 U355 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND23 U356 ( .A(n171), .B(n153), .Q(n151) );
  NAND26 U357 ( .A(n135), .B(n115), .Q(n113) );
  AOI212 U358 ( .A(n98), .B(n77), .C(n78), .Q(n429) );
  NOR22 U359 ( .A(n241), .B(n244), .Q(n239) );
  NOR24 U360 ( .A(B[8]), .B(n431), .Q(n244) );
  NOR24 U361 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NOR24 U362 ( .A(n113), .B(n151), .Q(n111) );
  NOR23 U363 ( .A(A[12]), .B(B[12]), .Q(n212) );
  AOI212 U364 ( .A(n443), .B(n55), .C(n56), .Q(n54) );
  NOR24 U365 ( .A(n88), .B(n79), .Q(n77) );
  AOI212 U366 ( .A(n443), .B(n97), .C(n420), .Q(n92) );
  NOR24 U367 ( .A(n439), .B(n435), .Q(n176) );
  BUF2 U368 ( .A(n205), .Q(n430) );
  INV4 U369 ( .A(n204), .Q(n440) );
  INV1 U370 ( .A(n429), .Q(n453) );
  OAI211 U371 ( .A(n70), .B(n416), .C(n71), .Q(n67) );
  INV2 U372 ( .A(n97), .Q(n458) );
  NAND28 U373 ( .A(n97), .B(n77), .Q(n6) );
  NOR23 U374 ( .A(n106), .B(n99), .Q(n97) );
  NOR23 U375 ( .A(n442), .B(n184), .Q(n182) );
  NOR23 U376 ( .A(n252), .B(n255), .Q(n250) );
  INV0 U377 ( .A(n145), .Q(n471) );
  NOR23 U378 ( .A(A[23]), .B(B[23]), .Q(n117) );
  NAND22 U379 ( .A(n111), .B(n66), .Q(n64) );
  INV3 U380 ( .A(n59), .Q(n450) );
  NOR23 U381 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR22 U382 ( .A(B[24]), .B(A[24]), .Q(n106) );
  BUF6 U383 ( .A(B[16]), .Q(n439) );
  BUF6 U384 ( .A(A[16]), .Q(n435) );
  NOR21 U385 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR22 U386 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR22 U387 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR23 U388 ( .A(n181), .B(n219), .Q(n179) );
  INV3 U389 ( .A(n244), .Q(n501) );
  AOI211 U390 ( .A(n472), .B(n135), .C(n436), .Q(n130) );
  NAND24 U391 ( .A(n423), .B(n65), .Q(n63) );
  BUF6 U392 ( .A(A[8]), .Q(n431) );
  BUF15 U393 ( .A(n178), .Q(n444) );
  NAND22 U394 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND21 U395 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND22 U396 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND22 U397 ( .A(B[19]), .B(A[19]), .Q(n156) );
  NAND22 U398 ( .A(B[25]), .B(A[25]), .Q(n100) );
  BUF2 U399 ( .A(n163), .Q(n433) );
  NOR24 U400 ( .A(B[19]), .B(A[19]), .Q(n432) );
  NOR24 U401 ( .A(n70), .B(n6), .Q(n66) );
  NAND22 U402 ( .A(B[17]), .B(A[17]), .Q(n174) );
  INV0 U404 ( .A(n126), .Q(n466) );
  INV0 U405 ( .A(n99), .Q(n457) );
  NAND24 U406 ( .A(n435), .B(n439), .Q(n177) );
  NOR24 U407 ( .A(n432), .B(n162), .Q(n153) );
  OAI212 U408 ( .A(n126), .B(n467), .C(n127), .Q(n123) );
  NAND21 U409 ( .A(n478), .B(n203), .Q(n197) );
  AOI210 U410 ( .A(n480), .B(n203), .C(n437), .Q(n198) );
  CLKIN3 U411 ( .A(n212), .Q(n486) );
  NAND24 U412 ( .A(n419), .B(n80), .Q(n78) );
  NAND24 U413 ( .A(n461), .B(n454), .Q(n419) );
  INV0 U414 ( .A(n223), .Q(n477) );
  AOI211 U415 ( .A(n472), .B(n122), .C(n123), .Q(n121) );
  NAND21 U416 ( .A(n474), .B(n122), .Q(n120) );
  INV0 U417 ( .A(n241), .Q(n498) );
  INV3 U418 ( .A(n436), .Q(n467) );
  CLKIN0 U419 ( .A(n480), .Q(n434) );
  INV0 U420 ( .A(n155), .Q(n473) );
  NOR21 U421 ( .A(n126), .B(n469), .Q(n122) );
  INV6 U422 ( .A(n183), .Q(n441) );
  NOR22 U423 ( .A(n173), .B(n176), .Q(n171) );
  CLKIN0 U424 ( .A(n417), .Q(n488) );
  XOR21 U425 ( .A(n22), .B(n444), .Q(SUM[16]) );
  INV6 U426 ( .A(n444), .Q(n479) );
  INV0 U427 ( .A(n173), .Q(n489) );
  CLKIN0 U428 ( .A(n176), .Q(n491) );
  NAND20 U429 ( .A(n177), .B(n491), .Q(n22) );
  NOR23 U430 ( .A(A[18]), .B(B[18]), .Q(n162) );
  NAND22 U431 ( .A(B[18]), .B(A[18]), .Q(n163) );
  NOR23 U432 ( .A(n61), .B(n70), .Q(n59) );
  INV1 U433 ( .A(n61), .Q(n449) );
  AOI212 U434 ( .A(n443), .B(n44), .C(n45), .Q(n43) );
  CLKIN0 U435 ( .A(n433), .Q(n476) );
  INV0 U436 ( .A(n117), .Q(n464) );
  OAI211 U437 ( .A(n145), .B(n137), .C(n138), .Q(n436) );
  OAI212 U438 ( .A(n219), .B(n495), .C(n434), .Q(n214) );
  NOR23 U439 ( .A(n205), .B(n212), .Q(n203) );
  NOR24 U440 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND22 U441 ( .A(B[14]), .B(A[14]), .Q(n195) );
  NOR21 U442 ( .A(n194), .B(n482), .Q(n190) );
  OAI211 U443 ( .A(n194), .B(n483), .C(n195), .Q(n191) );
  NOR22 U444 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NOR24 U445 ( .A(n117), .B(n126), .Q(n115) );
  NAND21 U446 ( .A(B[27]), .B(A[27]), .Q(n80) );
  CLKIN3 U447 ( .A(n106), .Q(n460) );
  NAND21 U448 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND22 U449 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND21 U450 ( .A(n446), .B(n51), .Q(n8) );
  AOI211 U451 ( .A(n480), .B(n190), .C(n191), .Q(n189) );
  OAI210 U452 ( .A(n177), .B(n173), .C(n174), .Q(n417) );
  XNR22 U453 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U454 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U455 ( .A(n15), .B(n119), .Q(SUM[23]) );
  XNR22 U456 ( .A(n20), .B(n164), .Q(SUM[18]) );
  XNR22 U457 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U458 ( .A(n475), .B(n433), .Q(n20) );
  INV0 U459 ( .A(n231), .Q(n493) );
  NOR24 U460 ( .A(B[9]), .B(A[9]), .Q(n241) );
  INV2 U461 ( .A(n88), .Q(n462) );
  NOR22 U462 ( .A(n88), .B(n458), .Q(n84) );
  NAND23 U463 ( .A(n59), .B(n446), .Q(n46) );
  AOI212 U464 ( .A(n60), .B(n446), .C(n447), .Q(n47) );
  INV2 U465 ( .A(n220), .Q(n480) );
  NAND24 U466 ( .A(n452), .B(n479), .Q(n423) );
  INV1 U467 ( .A(n230), .Q(n492) );
  NOR23 U468 ( .A(A[7]), .B(B[7]), .Q(n252) );
  CLKIN6 U469 ( .A(n79), .Q(n454) );
  NOR24 U470 ( .A(A[27]), .B(B[27]), .Q(n79) );
  NOR24 U471 ( .A(B[29]), .B(A[29]), .Q(n61) );
  AOI212 U472 ( .A(n443), .B(n84), .C(n85), .Q(n83) );
  AOI212 U473 ( .A(n443), .B(n455), .C(n453), .Q(n74) );
  INV2 U474 ( .A(n443), .Q(n463) );
  INV2 U475 ( .A(n144), .Q(n470) );
  INV2 U476 ( .A(n437), .Q(n483) );
  OAI211 U477 ( .A(n188), .B(n495), .C(n189), .Q(n187) );
  AOI212 U478 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U479 ( .A(n137), .B(n145), .C(n138), .Q(n136) );
  NOR24 U480 ( .A(n137), .B(n144), .Q(n135) );
  NOR24 U481 ( .A(B[21]), .B(A[21]), .Q(n137) );
  OAI212 U482 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  CLKIN0 U483 ( .A(n107), .Q(n459) );
  NAND21 U484 ( .A(n460), .B(n107), .Q(n14) );
  OAI211 U485 ( .A(n107), .B(n99), .C(n100), .Q(n420) );
  INV1 U486 ( .A(n162), .Q(n475) );
  AOI211 U487 ( .A(n472), .B(n470), .C(n471), .Q(n141) );
  INV2 U488 ( .A(n152), .Q(n472) );
  XNR22 U489 ( .A(n16), .B(n128), .Q(SUM[22]) );
  BUF15 U490 ( .A(n112), .Q(n443) );
  CLKIN1 U492 ( .A(n472), .Q(n438) );
  AOI212 U493 ( .A(n443), .B(n460), .C(n459), .Q(n103) );
  AOI210 U495 ( .A(n417), .B(n475), .C(n476), .Q(n159) );
  XNR22 U496 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR22 U497 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NOR24 U498 ( .A(B[19]), .B(A[19]), .Q(n155) );
  XNR22 U499 ( .A(n7), .B(n41), .Q(SUM[31]) );
  INV0 U500 ( .A(n255), .Q(n502) );
  OAI210 U501 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  XNR22 U502 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U503 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U504 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XNR22 U505 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NOR24 U506 ( .A(n440), .B(n441), .Q(n442) );
  NAND23 U507 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U508 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND22 U509 ( .A(n431), .B(B[8]), .Q(n245) );
  OAI212 U510 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NAND22 U511 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND21 U512 ( .A(n470), .B(n145), .Q(n18) );
  NAND21 U513 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV0 U514 ( .A(n185), .Q(n484) );
  OAI212 U515 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  NAND21 U516 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NOR24 U517 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND24 U518 ( .A(A[26]), .B(B[26]), .Q(n89) );
  OAI212 U519 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI210 U520 ( .A(n213), .B(n205), .C(n206), .Q(n437) );
  NOR24 U521 ( .A(A[17]), .B(B[17]), .Q(n173) );
  NOR24 U522 ( .A(A[13]), .B(B[13]), .Q(n205) );
  XNR22 U523 ( .A(n18), .B(n146), .Q(SUM[20]) );
  OAI212 U524 ( .A(n151), .B(n444), .C(n438), .Q(n146) );
  NAND24 U525 ( .A(n203), .B(n183), .Q(n181) );
  NOR24 U526 ( .A(n223), .B(n230), .Q(n221) );
  XNR22 U527 ( .A(n21), .B(n175), .Q(SUM[17]) );
  OAI212 U528 ( .A(n176), .B(n444), .C(n177), .Q(n175) );
  INV2 U529 ( .A(n70), .Q(n451) );
  NAND22 U530 ( .A(n481), .B(n206), .Q(n25) );
  NAND22 U531 ( .A(B[13]), .B(A[13]), .Q(n206) );
  NOR24 U532 ( .A(A[25]), .B(B[25]), .Q(n99) );
  INV4 U533 ( .A(n6), .Q(n455) );
  NOR22 U534 ( .A(n450), .B(n6), .Q(n55) );
  INV2 U535 ( .A(n135), .Q(n469) );
  NAND21 U536 ( .A(n474), .B(n135), .Q(n129) );
  AOI212 U537 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NOR22 U538 ( .A(n46), .B(n6), .Q(n44) );
  OAI212 U539 ( .A(n152), .B(n113), .C(n114), .Q(n112) );
  NAND24 U540 ( .A(n239), .B(n221), .Q(n219) );
  NOR24 U541 ( .A(A[22]), .B(B[22]), .Q(n126) );
  INV4 U542 ( .A(n247), .Q(n495) );
  OAI211 U543 ( .A(n450), .B(n429), .C(n448), .Q(n56) );
  OAI211 U544 ( .A(n46), .B(n416), .C(n47), .Q(n45) );
  AOI212 U545 ( .A(n443), .B(n66), .C(n67), .Q(n65) );
  OAI212 U546 ( .A(n444), .B(n91), .C(n92), .Q(n90) );
  NOR22 U547 ( .A(B[20]), .B(A[20]), .Q(n144) );
  OAI211 U548 ( .A(n244), .B(n495), .C(n245), .Q(n243) );
  AOI212 U549 ( .A(n98), .B(n77), .C(n78), .Q(n416) );
  INV0 U550 ( .A(n194), .Q(n485) );
  NOR24 U551 ( .A(n185), .B(n194), .Q(n183) );
  NAND21 U552 ( .A(B[7]), .B(A[7]), .Q(n253) );
  NOR23 U553 ( .A(B[15]), .B(A[15]), .Q(n185) );
  OAI211 U554 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  NAND22 U555 ( .A(A[6]), .B(B[6]), .Q(n256) );
  CLKIN0 U556 ( .A(n137), .Q(n468) );
  CLKIN0 U557 ( .A(n240), .Q(n500) );
  NAND22 U558 ( .A(n474), .B(n470), .Q(n140) );
  INV0 U559 ( .A(n171), .Q(n490) );
  NAND21 U560 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV0 U561 ( .A(n213), .Q(n487) );
  NAND20 U562 ( .A(n171), .B(n475), .Q(n158) );
  INV0 U563 ( .A(n430), .Q(n481) );
  INV0 U564 ( .A(n260), .Q(n497) );
  NOR20 U565 ( .A(n260), .B(n265), .Q(n258) );
  NAND21 U566 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U567 ( .A(n39), .Q(n445) );
  NAND21 U568 ( .A(n451), .B(n71), .Q(n10) );
  INV3 U569 ( .A(n219), .Q(n478) );
  INV3 U570 ( .A(n151), .Q(n474) );
  AOI211 U571 ( .A(n505), .B(n258), .C(n259), .Q(n257) );
  NAND22 U572 ( .A(n478), .B(n190), .Q(n188) );
  NAND20 U573 ( .A(n428), .B(n492), .Q(n226) );
  NAND22 U574 ( .A(n478), .B(n486), .Q(n208) );
  AOI210 U575 ( .A(n480), .B(n486), .C(n487), .Q(n209) );
  NAND22 U576 ( .A(n258), .B(n250), .Q(n248) );
  INV3 U577 ( .A(n420), .Q(n456) );
  INV3 U578 ( .A(n252), .Q(n503) );
  INV3 U579 ( .A(n64), .Q(n452) );
  INV3 U580 ( .A(n268), .Q(n505) );
  NAND22 U581 ( .A(A[10]), .B(B[10]), .Q(n231) );
  INV3 U582 ( .A(n51), .Q(n447) );
  CLKIN3 U583 ( .A(n89), .Q(n461) );
  NAND22 U584 ( .A(n497), .B(n261), .Q(n33) );
  INV3 U585 ( .A(n265), .Q(n496) );
  INV3 U586 ( .A(n274), .Q(n506) );
  NAND22 U587 ( .A(n504), .B(n272), .Q(n35) );
  INV3 U588 ( .A(n271), .Q(n504) );
  INV3 U589 ( .A(n266), .Q(n494) );
  AOI211 U590 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U591 ( .A(n271), .B(n274), .Q(n269) );
  INV3 U592 ( .A(n277), .Q(n508) );
  INV3 U593 ( .A(n278), .Q(n510) );
  NAND22 U594 ( .A(A[4]), .B(B[4]), .Q(n266) );
  INV3 U595 ( .A(n50), .Q(n446) );
  NOR21 U596 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U597 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U598 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U599 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U600 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U601 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND22 U602 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NOR21 U603 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U604 ( .A(A[0]), .B(B[0]), .Q(n281) );
  INV3 U605 ( .A(n280), .Q(n509) );
  NOR21 U606 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U607 ( .A(n462), .B(n89), .Q(n12) );
  NAND20 U608 ( .A(n449), .B(n62), .Q(n9) );
  NAND22 U609 ( .A(n445), .B(n40), .Q(n7) );
  NAND20 U610 ( .A(n454), .B(n80), .Q(n11) );
  NAND20 U611 ( .A(n489), .B(n174), .Q(n21) );
  XNR21 U612 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U613 ( .A(n486), .B(n213), .Q(n26) );
  XNR21 U614 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U615 ( .A(n484), .B(n186), .Q(n23) );
  XNR21 U616 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U617 ( .A(n477), .B(n224), .Q(n27) );
  XNR21 U618 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U619 ( .A(n498), .B(n242), .Q(n29) );
  XNR21 U620 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U621 ( .A(n485), .B(n195), .Q(n24) );
  XOR20 U622 ( .A(n30), .B(n495), .Q(SUM[8]) );
  NAND20 U623 ( .A(n245), .B(n501), .Q(n30) );
  XNR21 U624 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U625 ( .A(n492), .B(n231), .Q(n28) );
  XNR21 U626 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XNR21 U627 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U628 ( .A(n503), .B(n253), .Q(n31) );
  XOR21 U629 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND20 U630 ( .A(n502), .B(n256), .Q(n32) );
  NAND20 U631 ( .A(n464), .B(n118), .Q(n15) );
  NAND20 U632 ( .A(n156), .B(n473), .Q(n19) );
  NAND20 U633 ( .A(n466), .B(n127), .Q(n16) );
  XOR21 U634 ( .A(n36), .B(n508), .Q(SUM[2]) );
  NAND22 U635 ( .A(n506), .B(n275), .Q(n36) );
  XNR21 U636 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XOR21 U637 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U638 ( .A(n505), .B(n496), .C(n494), .Q(n262) );
  XNR21 U639 ( .A(n34), .B(n505), .Q(SUM[4]) );
  NAND22 U640 ( .A(n496), .B(n266), .Q(n34) );
  XOR21 U641 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U642 ( .A(n510), .B(n279), .Q(n37) );
  INV3 U643 ( .A(n38), .Q(SUM[0]) );
  NAND22 U644 ( .A(n509), .B(n281), .Q(n38) );
  NAND22 U645 ( .A(n111), .B(n460), .Q(n102) );
  NAND22 U646 ( .A(n111), .B(n84), .Q(n82) );
  NAND22 U647 ( .A(n111), .B(n55), .Q(n53) );
  NAND22 U648 ( .A(n111), .B(n455), .Q(n73) );
  NAND22 U649 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U650 ( .A(n111), .Q(n465) );
  AOI210 U651 ( .A(n240), .B(n492), .C(n493), .Q(n227) );
  NAND22 U652 ( .A(n468), .B(n138), .Q(n17) );
  NAND22 U653 ( .A(B[21]), .B(A[21]), .Q(n138) );
  OAI212 U654 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  INV2 U655 ( .A(n60), .Q(n448) );
endmodule


module adder_44 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_44_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_43_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n205, n206, n207, n208, n209, n212, n213,
         n214, n219, n220, n221, n222, n223, n224, n225, n226, n227, n230,
         n231, n232, n239, n240, n241, n242, n243, n244, n245, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n265, n266, n268, n269, n270, n271, n272, n273,
         n274, n275, n277, n278, n279, n280, n281, n420, n421, n422, n433,
         n434, n438, n439, n442, n443, n449, n450, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n603, n604, n605, n606, n607, n608;

  OAI212 U51 ( .A(n73), .B(n537), .C(n74), .Q(n72) );
  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U65 ( .A(n82), .B(n537), .C(n83), .Q(n81) );
  OAI212 U77 ( .A(n91), .B(n537), .C(n92), .Q(n90) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U91 ( .A(n102), .B(n537), .C(n103), .Q(n101) );
  OAI212 U101 ( .A(n554), .B(n537), .C(n552), .Q(n108) );
  OAI212 U115 ( .A(n120), .B(n537), .C(n121), .Q(n119) );
  OAI212 U127 ( .A(n129), .B(n537), .C(n130), .Q(n128) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n537), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U159 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U165 ( .A(n158), .B(n537), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n572), .B(n537), .C(n570), .Q(n164) );
  OAI212 U183 ( .A(n531), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U201 ( .A(n530), .B(n185), .C(n186), .Q(n184) );
  OAI212 U207 ( .A(n188), .B(n574), .C(n189), .Q(n187) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n266), .B(n534), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n604), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U411 ( .A(n213), .B(n205), .C(n206), .Q(n422) );
  OAI212 U500 ( .A(n176), .B(n537), .C(n531), .Q(n175) );
  OAI212 U442 ( .A(n42), .B(n537), .C(n43), .Q(n41) );
  CLKBU12 U349 ( .A(n195), .Q(n530) );
  NOR21 U350 ( .A(n61), .B(n70), .Q(n59) );
  NOR22 U351 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NAND22 U352 ( .A(A[11]), .B(B[11]), .Q(n224) );
  XNR22 U353 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NOR22 U354 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND21 U355 ( .A(A[14]), .B(B[14]), .Q(n195) );
  CLKIN4 U356 ( .A(n175), .Q(n559) );
  XOR21 U357 ( .A(n30), .B(n574), .Q(SUM[8]) );
  INV8 U358 ( .A(n247), .Q(n574) );
  BUF15 U359 ( .A(n178), .Q(n537) );
  NOR24 U360 ( .A(B[9]), .B(A[9]), .Q(n241) );
  OAI210 U361 ( .A(n126), .B(n567), .C(n127), .Q(n123) );
  NAND22 U362 ( .A(n175), .B(n21), .Q(n438) );
  CLKIN3 U363 ( .A(n203), .Q(n595) );
  NOR22 U364 ( .A(n173), .B(n176), .Q(n171) );
  NOR24 U365 ( .A(n155), .B(n162), .Q(n153) );
  NOR22 U366 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NAND24 U367 ( .A(n528), .B(n203), .Q(n181) );
  AOI211 U368 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR22 U369 ( .A(n79), .B(n88), .Q(n77) );
  NOR23 U370 ( .A(n113), .B(n151), .Q(n111) );
  INV3 U371 ( .A(n219), .Q(n578) );
  BUF8 U372 ( .A(n194), .Q(n532) );
  BUF8 U373 ( .A(n111), .Q(n535) );
  NOR21 U374 ( .A(n585), .B(n6), .Q(n55) );
  NAND23 U375 ( .A(n171), .B(n153), .Q(n151) );
  NAND24 U376 ( .A(n544), .B(n548), .Q(n443) );
  INV3 U377 ( .A(n565), .Q(n517) );
  NAND21 U378 ( .A(B[7]), .B(A[7]), .Q(n253) );
  NAND22 U379 ( .A(n157), .B(n19), .Q(n420) );
  NAND26 U380 ( .A(n558), .B(n562), .Q(n421) );
  INV2 U381 ( .A(n583), .Q(n518) );
  INV2 U382 ( .A(n240), .Q(n583) );
  CLKIN4 U383 ( .A(n157), .Q(n558) );
  INV2 U384 ( .A(n570), .Q(n519) );
  INV1 U385 ( .A(n172), .Q(n570) );
  NAND23 U386 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND20 U387 ( .A(n593), .B(n224), .Q(n27) );
  NOR24 U388 ( .A(B[11]), .B(A[11]), .Q(n223) );
  CLKIN4 U389 ( .A(n81), .Q(n543) );
  NAND21 U390 ( .A(A[13]), .B(B[13]), .Q(n206) );
  INV3 U391 ( .A(n185), .Q(n591) );
  NAND21 U392 ( .A(A[15]), .B(B[15]), .Q(n186) );
  INV2 U393 ( .A(n152), .Q(n565) );
  NAND20 U394 ( .A(n563), .B(n156), .Q(n19) );
  NAND22 U395 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NOR22 U396 ( .A(n252), .B(n255), .Q(n250) );
  NAND22 U397 ( .A(n101), .B(n13), .Q(n522) );
  NAND23 U398 ( .A(n520), .B(n521), .Q(n523) );
  NAND24 U399 ( .A(n522), .B(n523), .Q(SUM[25]) );
  CLKIN3 U400 ( .A(n101), .Q(n520) );
  INV3 U401 ( .A(n13), .Q(n521) );
  OAI211 U402 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI211 U403 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NAND21 U404 ( .A(n592), .B(n256), .Q(n32) );
  NAND21 U405 ( .A(A[24]), .B(B[24]), .Q(n107) );
  CLKIN0 U406 ( .A(n223), .Q(n593) );
  NOR24 U407 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR20 U408 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND22 U409 ( .A(n24), .B(n196), .Q(n526) );
  NAND26 U410 ( .A(n524), .B(n525), .Q(n527) );
  NAND28 U412 ( .A(n526), .B(n527), .Q(SUM[14]) );
  INV6 U413 ( .A(n24), .Q(n524) );
  CLKIN6 U414 ( .A(n196), .Q(n525) );
  NAND21 U415 ( .A(n557), .B(n530), .Q(n24) );
  INV0 U416 ( .A(n241), .Q(n588) );
  AOI212 U417 ( .A(n433), .B(n551), .C(n550), .Q(n103) );
  NAND22 U418 ( .A(n258), .B(n250), .Q(n248) );
  NOR20 U419 ( .A(B[4]), .B(A[4]), .Q(n265) );
  CLKIN4 U420 ( .A(n90), .Q(n548) );
  OAI212 U421 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  INV2 U422 ( .A(n205), .Q(n598) );
  NOR23 U423 ( .A(B[13]), .B(A[13]), .Q(n205) );
  OAI212 U424 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  NOR23 U425 ( .A(n185), .B(n532), .Q(n183) );
  NAND28 U426 ( .A(n438), .B(n439), .Q(SUM[17]) );
  NAND22 U427 ( .A(n577), .B(n231), .Q(n28) );
  NAND22 U428 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND21 U429 ( .A(A[26]), .B(B[26]), .Q(n89) );
  XOR22 U430 ( .A(n22), .B(n537), .Q(SUM[16]) );
  NOR23 U431 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR22 U432 ( .A(n532), .B(n595), .Q(n190) );
  CLKIN0 U433 ( .A(n532), .Q(n557) );
  NAND20 U434 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV6 U435 ( .A(n220), .Q(n579) );
  OAI211 U436 ( .A(n532), .B(n597), .C(n530), .Q(n191) );
  BUF4 U437 ( .A(n111), .Q(n536) );
  NOR23 U438 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR24 U439 ( .A(n185), .B(n532), .Q(n528) );
  NOR23 U440 ( .A(n223), .B(n230), .Q(n221) );
  NAND28 U441 ( .A(n442), .B(n443), .Q(SUM[26]) );
  CLKBU12 U443 ( .A(n177), .Q(n531) );
  NAND21 U444 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NOR23 U445 ( .A(n241), .B(n244), .Q(n239) );
  AOI211 U446 ( .A(n433), .B(n55), .C(n56), .Q(n54) );
  OAI211 U447 ( .A(n53), .B(n537), .C(n54), .Q(n52) );
  INV0 U448 ( .A(n252), .Q(n573) );
  AOI211 U449 ( .A(n565), .B(n135), .C(n136), .Q(n130) );
  NAND28 U450 ( .A(n449), .B(n450), .Q(SUM[27]) );
  NAND26 U451 ( .A(n543), .B(n539), .Q(n450) );
  NAND22 U452 ( .A(n81), .B(n11), .Q(n449) );
  AOI212 U453 ( .A(n433), .B(n84), .C(n85), .Q(n83) );
  OAI212 U454 ( .A(n113), .B(n152), .C(n114), .Q(n433) );
  INV1 U455 ( .A(n230), .Q(n577) );
  NOR22 U456 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND28 U457 ( .A(n135), .B(n115), .Q(n113) );
  NOR24 U458 ( .A(n117), .B(n126), .Q(n115) );
  XNR22 U459 ( .A(n10), .B(n72), .Q(SUM[28]) );
  OAI212 U460 ( .A(n197), .B(n574), .C(n198), .Q(n196) );
  XNR22 U461 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NOR21 U462 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND26 U463 ( .A(n559), .B(n589), .Q(n439) );
  NAND21 U464 ( .A(A[22]), .B(B[22]), .Q(n127) );
  AOI211 U465 ( .A(n112), .B(n541), .C(n542), .Q(n74) );
  INV1 U466 ( .A(n5), .Q(n542) );
  INV1 U467 ( .A(n579), .Q(n529) );
  NAND28 U468 ( .A(n420), .B(n421), .Q(SUM[19]) );
  NAND23 U469 ( .A(n239), .B(n221), .Q(n219) );
  NAND20 U470 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NOR22 U471 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND20 U472 ( .A(A[19]), .B(B[19]), .Q(n156) );
  OAI212 U473 ( .A(n151), .B(n537), .C(n517), .Q(n146) );
  NOR23 U474 ( .A(n181), .B(n219), .Q(n179) );
  XNR22 U475 ( .A(n20), .B(n164), .Q(SUM[18]) );
  OAI212 U476 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NOR22 U477 ( .A(B[27]), .B(A[27]), .Q(n79) );
  XNR22 U478 ( .A(n17), .B(n139), .Q(SUM[21]) );
  OAI212 U479 ( .A(n208), .B(n574), .C(n209), .Q(n207) );
  AOI211 U480 ( .A(n579), .B(n594), .C(n596), .Q(n209) );
  NOR23 U481 ( .A(n99), .B(n106), .Q(n97) );
  INV0 U482 ( .A(n99), .Q(n546) );
  OAI211 U483 ( .A(n64), .B(n537), .C(n65), .Q(n63) );
  AOI211 U484 ( .A(n112), .B(n66), .C(n67), .Q(n65) );
  NOR22 U485 ( .A(B[16]), .B(A[16]), .Q(n176) );
  INV2 U486 ( .A(n126), .Q(n556) );
  NOR22 U487 ( .A(B[22]), .B(A[22]), .Q(n126) );
  XNR22 U488 ( .A(n29), .B(n243), .Q(SUM[9]) );
  XNR22 U489 ( .A(n26), .B(n214), .Q(SUM[12]) );
  AOI212 U490 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  XNR22 U491 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U492 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND20 U493 ( .A(n545), .B(n89), .Q(n12) );
  OAI211 U494 ( .A(n88), .B(n549), .C(n89), .Q(n85) );
  OAI211 U495 ( .A(n585), .B(n5), .C(n586), .Q(n56) );
  OAI210 U496 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  NOR23 U497 ( .A(n137), .B(n144), .Q(n135) );
  NOR21 U498 ( .A(B[20]), .B(A[20]), .Q(n144) );
  INV2 U499 ( .A(n212), .Q(n594) );
  INV0 U501 ( .A(n176), .Q(n571) );
  XNR22 U502 ( .A(n23), .B(n187), .Q(SUM[15]) );
  XNR22 U503 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NAND21 U504 ( .A(n594), .B(n213), .Q(n26) );
  CLKIN2 U505 ( .A(n213), .Q(n596) );
  NAND22 U506 ( .A(A[12]), .B(B[12]), .Q(n213) );
  INV2 U507 ( .A(n422), .Q(n597) );
  NOR22 U508 ( .A(B[23]), .B(A[23]), .Q(n117) );
  OAI211 U509 ( .A(n219), .B(n574), .C(n529), .Q(n214) );
  AOI212 U510 ( .A(n221), .B(n240), .C(n222), .Q(n220) );
  XNR22 U511 ( .A(n15), .B(n119), .Q(SUM[23]) );
  INV2 U512 ( .A(n151), .Q(n564) );
  OAI211 U513 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND22 U514 ( .A(n535), .B(n55), .Q(n53) );
  XNR22 U515 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NOR23 U516 ( .A(n205), .B(n212), .Q(n203) );
  NOR24 U517 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND22 U518 ( .A(n535), .B(n66), .Q(n64) );
  AOI212 U519 ( .A(n183), .B(n422), .C(n184), .Q(n182) );
  XNR22 U520 ( .A(n18), .B(n146), .Q(SUM[20]) );
  INV0 U521 ( .A(n117), .Q(n553) );
  OAI211 U522 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NAND21 U523 ( .A(A[18]), .B(B[18]), .Q(n163) );
  OAI211 U524 ( .A(n582), .B(n574), .C(n583), .Q(n232) );
  OAI211 U525 ( .A(n226), .B(n574), .C(n227), .Q(n225) );
  OAI211 U526 ( .A(n244), .B(n574), .C(n245), .Q(n243) );
  XNR22 U527 ( .A(n25), .B(n207), .Q(SUM[13]) );
  INV2 U528 ( .A(n6), .Q(n541) );
  CLKIN1 U529 ( .A(n98), .Q(n549) );
  NAND21 U530 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U531 ( .A(n578), .B(n190), .Q(n188) );
  NAND21 U532 ( .A(n578), .B(n203), .Q(n197) );
  CLKIN1 U533 ( .A(n536), .Q(n554) );
  NAND20 U534 ( .A(n540), .B(n80), .Q(n11) );
  CLKIN3 U535 ( .A(n534), .Q(n601) );
  NAND21 U536 ( .A(n536), .B(n541), .Q(n73) );
  NAND22 U537 ( .A(n564), .B(n555), .Q(n120) );
  NAND20 U538 ( .A(n171), .B(n576), .Q(n158) );
  INV0 U539 ( .A(n163), .Q(n575) );
  NAND22 U540 ( .A(n564), .B(n135), .Q(n129) );
  NAND21 U541 ( .A(n587), .B(n71), .Q(n10) );
  NAND22 U542 ( .A(n584), .B(n62), .Q(n9) );
  INV0 U543 ( .A(n61), .Q(n584) );
  NOR20 U544 ( .A(B[20]), .B(A[20]), .Q(n533) );
  AOI210 U545 ( .A(n579), .B(n203), .C(n422), .Q(n198) );
  NAND21 U546 ( .A(n568), .B(n145), .Q(n18) );
  INV2 U547 ( .A(n21), .Q(n589) );
  NAND21 U548 ( .A(n576), .B(n163), .Q(n20) );
  NAND20 U549 ( .A(n556), .B(n135), .Q(n434) );
  INV0 U550 ( .A(n244), .Q(n581) );
  NAND20 U551 ( .A(n556), .B(n127), .Q(n16) );
  INV0 U552 ( .A(n70), .Q(n587) );
  NAND20 U553 ( .A(n551), .B(n107), .Q(n14) );
  AOI210 U554 ( .A(n60), .B(n561), .C(n560), .Q(n47) );
  NOR20 U555 ( .A(n534), .B(n265), .Q(n258) );
  NAND20 U556 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U557 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U558 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND20 U559 ( .A(n536), .B(n44), .Q(n42) );
  NAND22 U560 ( .A(n239), .B(n577), .Q(n226) );
  NAND22 U561 ( .A(n578), .B(n594), .Q(n208) );
  NAND22 U562 ( .A(n564), .B(n568), .Q(n140) );
  INV3 U563 ( .A(n239), .Q(n582) );
  XNR21 U564 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U565 ( .A(n573), .B(n253), .Q(n31) );
  NAND20 U566 ( .A(n581), .B(n245), .Q(n30) );
  NAND20 U567 ( .A(n588), .B(n242), .Q(n29) );
  XOR21 U568 ( .A(n32), .B(n257), .Q(SUM[6]) );
  INV2 U569 ( .A(n255), .Q(n592) );
  NAND20 U570 ( .A(n598), .B(n206), .Q(n25) );
  NAND20 U571 ( .A(n591), .B(n186), .Q(n23) );
  NAND22 U572 ( .A(n97), .B(n77), .Q(n6) );
  INV3 U573 ( .A(n145), .Q(n569) );
  NOR20 U574 ( .A(n46), .B(n6), .Q(n44) );
  NAND22 U575 ( .A(n535), .B(n97), .Q(n91) );
  AOI211 U576 ( .A(n112), .B(n97), .C(n98), .Q(n92) );
  AOI211 U577 ( .A(n579), .B(n190), .C(n191), .Q(n189) );
  NAND20 U578 ( .A(n590), .B(n174), .Q(n21) );
  INV3 U579 ( .A(n173), .Q(n590) );
  INV3 U580 ( .A(n60), .Q(n586) );
  AOI210 U581 ( .A(n518), .B(n577), .C(n580), .Q(n227) );
  INV0 U582 ( .A(n231), .Q(n580) );
  INV3 U583 ( .A(n11), .Q(n539) );
  NAND22 U584 ( .A(n12), .B(n90), .Q(n442) );
  INV3 U585 ( .A(n12), .Q(n544) );
  INV3 U586 ( .A(n533), .Q(n568) );
  INV3 U587 ( .A(n19), .Q(n562) );
  INV3 U588 ( .A(n162), .Q(n576) );
  INV3 U589 ( .A(n171), .Q(n572) );
  INV3 U590 ( .A(n59), .Q(n585) );
  NAND22 U591 ( .A(n536), .B(n551), .Q(n102) );
  INV3 U592 ( .A(n97), .Q(n547) );
  INV3 U593 ( .A(n434), .Q(n555) );
  AOI211 U594 ( .A(n605), .B(n258), .C(n259), .Q(n257) );
  INV3 U595 ( .A(n268), .Q(n605) );
  INV3 U596 ( .A(n277), .Q(n604) );
  NAND22 U597 ( .A(n571), .B(n531), .Q(n22) );
  NOR21 U598 ( .A(n70), .B(n6), .Q(n66) );
  NAND20 U599 ( .A(n546), .B(n100), .Q(n13) );
  XNR21 U600 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND22 U601 ( .A(n561), .B(n51), .Q(n8) );
  XNR21 U602 ( .A(n34), .B(n605), .Q(SUM[4]) );
  NAND22 U603 ( .A(n599), .B(n266), .Q(n34) );
  NAND20 U604 ( .A(n566), .B(n138), .Q(n17) );
  INV0 U605 ( .A(n137), .Q(n566) );
  NAND22 U606 ( .A(n553), .B(n118), .Q(n15) );
  CLKIN2 U607 ( .A(n106), .Q(n551) );
  INV3 U608 ( .A(n79), .Q(n540) );
  INV0 U609 ( .A(n88), .Q(n545) );
  NAND21 U610 ( .A(n535), .B(n84), .Q(n82) );
  NOR21 U611 ( .A(n88), .B(n547), .Q(n84) );
  INV0 U612 ( .A(n155), .Q(n563) );
  INV3 U613 ( .A(n107), .Q(n550) );
  INV3 U614 ( .A(n265), .Q(n599) );
  AOI210 U615 ( .A(n433), .B(n44), .C(n45), .Q(n43) );
  INV3 U616 ( .A(n51), .Q(n560) );
  AOI211 U617 ( .A(n565), .B(n555), .C(n123), .Q(n121) );
  INV0 U618 ( .A(n136), .Q(n567) );
  NAND21 U619 ( .A(n59), .B(n561), .Q(n46) );
  XOR21 U620 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U621 ( .A(n605), .B(n599), .C(n600), .Q(n262) );
  NAND22 U622 ( .A(n601), .B(n261), .Q(n33) );
  INV3 U623 ( .A(n266), .Q(n600) );
  AOI211 U624 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U625 ( .A(n271), .B(n274), .Q(n269) );
  XOR21 U626 ( .A(n36), .B(n604), .Q(SUM[2]) );
  NAND22 U627 ( .A(n607), .B(n275), .Q(n36) );
  INV3 U628 ( .A(n274), .Q(n607) );
  XOR21 U629 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U630 ( .A(n606), .B(n279), .Q(n37) );
  INV3 U631 ( .A(n278), .Q(n606) );
  XNR21 U632 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U633 ( .A(n608), .B(n272), .Q(n35) );
  INV3 U634 ( .A(n271), .Q(n608) );
  NAND20 U635 ( .A(A[28]), .B(B[28]), .Q(n71) );
  XNR21 U636 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U637 ( .A(n538), .B(n40), .Q(n7) );
  NAND20 U638 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND20 U639 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV3 U640 ( .A(n50), .Q(n561) );
  BUF2 U641 ( .A(n260), .Q(n534) );
  INV3 U642 ( .A(n39), .Q(n538) );
  NOR20 U643 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U644 ( .A(n38), .Q(SUM[0]) );
  NAND22 U645 ( .A(n603), .B(n281), .Q(n38) );
  INV3 U646 ( .A(n280), .Q(n603) );
  NOR20 U647 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NOR20 U648 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR20 U649 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND20 U650 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U651 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NOR20 U652 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND20 U653 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U654 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND21 U655 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NOR20 U656 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND22 U657 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND22 U658 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NOR21 U659 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR22 U660 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR22 U661 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR20 U662 ( .A(B[5]), .B(A[5]), .Q(n260) );
  AOI210 U663 ( .A(n519), .B(n576), .C(n575), .Q(n159) );
  INV1 U664 ( .A(n112), .Q(n552) );
  AOI211 U665 ( .A(n565), .B(n568), .C(n569), .Q(n141) );
  NOR22 U666 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR22 U667 ( .A(B[21]), .B(A[21]), .Q(n137) );
endmodule


module adder_43 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_43_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_42_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n418, n419, n423,
         n426, n427, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n518, n519, n520;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U59 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U77 ( .A(n91), .B(n450), .C(n92), .Q(n90) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U91 ( .A(n102), .B(n450), .C(n103), .Q(n101) );
  OAI212 U101 ( .A(n468), .B(n450), .C(n466), .Q(n108) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U127 ( .A(n129), .B(n450), .C(n130), .Q(n128) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n450), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n450), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n492), .B(n450), .C(n493), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n221), .B(n240), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n502), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n515), .B(n502), .C(n513), .Q(n232) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  AOI212 U290 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U329 ( .A(n274), .B(n519), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U352 ( .A(n73), .B(n450), .C(n74), .Q(n72) );
  OAI212 U507 ( .A(n53), .B(n442), .C(n54), .Q(n52) );
  OAI211 U349 ( .A(n456), .B(n5), .C(n454), .Q(n56) );
  XNR22 U350 ( .A(n28), .B(n232), .Q(SUM[10]) );
  CLKIN4 U351 ( .A(n157), .Q(n481) );
  NOR24 U353 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND23 U354 ( .A(A[16]), .B(B[16]), .Q(n177) );
  XNR22 U355 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NOR22 U356 ( .A(n70), .B(n6), .Q(n66) );
  AOI212 U357 ( .A(n97), .B(n434), .C(n98), .Q(n92) );
  INV4 U358 ( .A(n502), .Q(n439) );
  NOR23 U359 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR24 U360 ( .A(n260), .B(n265), .Q(n258) );
  XNR22 U361 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NOR23 U362 ( .A(n155), .B(n162), .Q(n153) );
  INV2 U363 ( .A(n230), .Q(n488) );
  NOR24 U364 ( .A(n252), .B(n255), .Q(n250) );
  NOR23 U365 ( .A(n173), .B(n176), .Q(n171) );
  NOR22 U366 ( .A(B[27]), .B(A[27]), .Q(n79) );
  INV1 U367 ( .A(n162), .Q(n482) );
  NAND21 U368 ( .A(n480), .B(n423), .Q(n140) );
  INV6 U369 ( .A(n423), .Q(n473) );
  AOI211 U370 ( .A(n478), .B(n423), .C(n475), .Q(n141) );
  NAND28 U371 ( .A(n476), .B(n474), .Q(n423) );
  OAI211 U372 ( .A(n126), .B(n470), .C(n127), .Q(n123) );
  NAND26 U373 ( .A(n135), .B(n115), .Q(n113) );
  AOI212 U374 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NOR23 U375 ( .A(n117), .B(n126), .Q(n115) );
  NAND24 U376 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND24 U377 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND24 U378 ( .A(n503), .B(n505), .Q(n430) );
  NAND22 U379 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND24 U380 ( .A(n438), .B(n439), .Q(n440) );
  NAND22 U381 ( .A(n97), .B(n77), .Q(n6) );
  NOR22 U382 ( .A(B[23]), .B(A[23]), .Q(n117) );
  INV3 U383 ( .A(n90), .Q(n463) );
  NOR21 U384 ( .A(B[29]), .B(A[29]), .Q(n61) );
  AOI211 U385 ( .A(n435), .B(n461), .C(n464), .Q(n103) );
  NOR21 U386 ( .A(n456), .B(n6), .Q(n55) );
  AOI211 U387 ( .A(n435), .B(n84), .C(n85), .Q(n83) );
  NOR22 U388 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR22 U389 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND22 U390 ( .A(n171), .B(n153), .Q(n151) );
  NOR22 U391 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR23 U392 ( .A(n113), .B(n151), .Q(n111) );
  NAND26 U393 ( .A(n481), .B(n477), .Q(n419) );
  INV3 U394 ( .A(n22), .Q(n448) );
  INV3 U395 ( .A(n484), .Q(n449) );
  INV3 U396 ( .A(n25), .Q(n447) );
  INV6 U397 ( .A(n112), .Q(n433) );
  INV3 U398 ( .A(n433), .Q(n434) );
  INV6 U399 ( .A(n433), .Q(n435) );
  INV1 U400 ( .A(n135), .Q(n472) );
  NOR24 U401 ( .A(B[13]), .B(A[13]), .Q(n205) );
  OAI211 U402 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI211 U403 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  CLKBU2 U404 ( .A(n259), .Q(n436) );
  INV2 U405 ( .A(n513), .Q(n437) );
  INV2 U406 ( .A(n240), .Q(n513) );
  INV1 U407 ( .A(n435), .Q(n466) );
  NOR23 U408 ( .A(B[19]), .B(A[19]), .Q(n155) );
  INV1 U409 ( .A(n98), .Q(n465) );
  OAI212 U410 ( .A(n64), .B(n450), .C(n65), .Q(n63) );
  NOR24 U411 ( .A(n223), .B(n230), .Q(n221) );
  NOR23 U412 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NAND20 U413 ( .A(n461), .B(n107), .Q(n14) );
  CLKIN3 U414 ( .A(n107), .Q(n464) );
  NAND20 U415 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NOR24 U416 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NOR22 U417 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV2 U418 ( .A(n204), .Q(n498) );
  NOR23 U419 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND22 U420 ( .A(A[18]), .B(B[18]), .Q(n163) );
  INV3 U421 ( .A(n220), .Q(n484) );
  NOR22 U422 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NAND22 U423 ( .A(n111), .B(n84), .Q(n82) );
  NAND21 U424 ( .A(n488), .B(n231), .Q(n28) );
  NAND28 U425 ( .A(n445), .B(n446), .Q(SUM[17]) );
  NAND21 U426 ( .A(A[24]), .B(B[24]), .Q(n107) );
  INV0 U427 ( .A(n223), .Q(n485) );
  NOR22 U428 ( .A(B[10]), .B(A[10]), .Q(n230) );
  CLKIN3 U429 ( .A(n175), .Q(n443) );
  NAND26 U430 ( .A(n440), .B(n209), .Q(n207) );
  INV3 U431 ( .A(n208), .Q(n438) );
  NAND23 U432 ( .A(n486), .B(n500), .Q(n208) );
  INV15 U433 ( .A(n247), .Q(n502) );
  OAI212 U434 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI211 U435 ( .A(n194), .B(n498), .C(n195), .Q(n191) );
  CLKIN3 U436 ( .A(n79), .Q(n458) );
  NOR23 U437 ( .A(B[6]), .B(A[6]), .Q(n255) );
  INV2 U438 ( .A(n152), .Q(n478) );
  CLKIN2 U439 ( .A(n450), .Q(n441) );
  INV3 U440 ( .A(n441), .Q(n442) );
  NAND22 U441 ( .A(n175), .B(n21), .Q(n445) );
  NAND24 U442 ( .A(n443), .B(n444), .Q(n446) );
  INV3 U443 ( .A(n21), .Q(n444) );
  NAND20 U444 ( .A(n482), .B(n163), .Q(n20) );
  INV2 U445 ( .A(n163), .Q(n483) );
  NAND21 U446 ( .A(n111), .B(n461), .Q(n102) );
  INV1 U447 ( .A(n106), .Q(n461) );
  NAND24 U448 ( .A(n239), .B(n221), .Q(n219) );
  NOR23 U449 ( .A(n181), .B(n219), .Q(n179) );
  NOR23 U450 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND22 U451 ( .A(n500), .B(n213), .Q(n26) );
  NAND22 U452 ( .A(A[12]), .B(B[12]), .Q(n213) );
  INV1 U453 ( .A(n241), .Q(n516) );
  XNR22 U454 ( .A(n448), .B(n450), .Q(SUM[16]) );
  XOR22 U455 ( .A(n447), .B(n207), .Q(SUM[13]) );
  OAI210 U456 ( .A(n42), .B(n442), .C(n43), .Q(n41) );
  NAND21 U457 ( .A(A[21]), .B(B[21]), .Q(n138) );
  AOI212 U458 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND24 U459 ( .A(n258), .B(n250), .Q(n248) );
  OAI211 U460 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  XNR22 U461 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NAND24 U462 ( .A(n203), .B(n183), .Q(n181) );
  NOR23 U463 ( .A(n185), .B(n194), .Q(n183) );
  NAND22 U464 ( .A(A[6]), .B(B[6]), .Q(n256) );
  OAI212 U465 ( .A(n244), .B(n502), .C(n245), .Q(n243) );
  NOR24 U466 ( .A(n205), .B(n212), .Q(n203) );
  NOR23 U467 ( .A(B[14]), .B(A[14]), .Q(n194) );
  XNR21 U468 ( .A(n34), .B(n505), .Q(SUM[4]) );
  AOI212 U469 ( .A(n505), .B(n258), .C(n436), .Q(n257) );
  NOR22 U470 ( .A(B[26]), .B(A[26]), .Q(n88) );
  OAI211 U471 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  INV0 U472 ( .A(n213), .Q(n499) );
  INV6 U473 ( .A(n248), .Q(n503) );
  NAND21 U474 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U475 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND22 U476 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND26 U477 ( .A(n489), .B(n463), .Q(n427) );
  NAND28 U478 ( .A(n426), .B(n427), .Q(SUM[26]) );
  BUF15 U479 ( .A(n178), .Q(n450) );
  NOR24 U480 ( .A(B[7]), .B(A[7]), .Q(n252) );
  INV6 U481 ( .A(A[20]), .Q(n474) );
  AOI211 U482 ( .A(n435), .B(n66), .C(n67), .Q(n65) );
  NAND21 U483 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NAND21 U484 ( .A(A[22]), .B(B[22]), .Q(n127) );
  AOI211 U485 ( .A(n435), .B(n55), .C(n56), .Q(n54) );
  OAI212 U486 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  AOI211 U487 ( .A(n478), .B(n122), .C(n123), .Q(n121) );
  NAND28 U488 ( .A(n418), .B(n419), .Q(SUM[19]) );
  NAND22 U489 ( .A(n157), .B(n19), .Q(n418) );
  NAND28 U490 ( .A(n430), .B(n249), .Q(n247) );
  OAI212 U491 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  AOI212 U492 ( .A(n484), .B(n500), .C(n499), .Q(n209) );
  XNR22 U493 ( .A(n9), .B(n63), .Q(SUM[29]) );
  CLKIN2 U494 ( .A(n203), .Q(n497) );
  INV2 U495 ( .A(B[20]), .Q(n476) );
  NAND24 U496 ( .A(A[7]), .B(B[7]), .Q(n253) );
  OAI212 U497 ( .A(n197), .B(n502), .C(n198), .Q(n196) );
  NAND21 U498 ( .A(A[11]), .B(B[11]), .Q(n224) );
  OAI212 U499 ( .A(n120), .B(n450), .C(n121), .Q(n119) );
  OAI212 U500 ( .A(n151), .B(n450), .C(n152), .Q(n146) );
  XNR22 U501 ( .A(n14), .B(n108), .Q(SUM[24]) );
  OAI212 U502 ( .A(n176), .B(n450), .C(n177), .Q(n175) );
  OAI212 U503 ( .A(n188), .B(n502), .C(n189), .Q(n187) );
  NAND22 U504 ( .A(n486), .B(n190), .Q(n188) );
  INV6 U505 ( .A(n268), .Q(n505) );
  NAND20 U506 ( .A(n495), .B(n174), .Q(n21) );
  XNR22 U508 ( .A(n8), .B(n52), .Q(SUM[30]) );
  OAI212 U509 ( .A(n219), .B(n502), .C(n449), .Q(n214) );
  AOI211 U510 ( .A(n484), .B(n190), .C(n191), .Q(n189) );
  OAI212 U511 ( .A(n450), .B(n82), .C(n83), .Q(n81) );
  OAI212 U512 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  AOI212 U513 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR22 U514 ( .A(n271), .B(n274), .Q(n269) );
  NAND20 U515 ( .A(n469), .B(n127), .Q(n16) );
  OAI211 U516 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  AOI211 U517 ( .A(n484), .B(n203), .C(n204), .Q(n198) );
  XNR22 U518 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND22 U519 ( .A(n111), .B(n66), .Q(n64) );
  XNR22 U520 ( .A(n20), .B(n164), .Q(SUM[18]) );
  XNR22 U521 ( .A(n29), .B(n243), .Q(SUM[9]) );
  XNR22 U522 ( .A(n13), .B(n101), .Q(SUM[25]) );
  AOI211 U523 ( .A(n435), .B(n459), .C(n460), .Q(n74) );
  XNR22 U524 ( .A(n26), .B(n214), .Q(SUM[12]) );
  XNR22 U525 ( .A(n15), .B(n119), .Q(SUM[23]) );
  INV3 U526 ( .A(n151), .Q(n480) );
  XNR22 U527 ( .A(n81), .B(n11), .Q(SUM[27]) );
  NAND21 U528 ( .A(n111), .B(n459), .Q(n73) );
  NOR23 U529 ( .A(B[8]), .B(A[8]), .Q(n244) );
  XNR22 U530 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NOR22 U531 ( .A(n79), .B(n88), .Q(n77) );
  NOR24 U532 ( .A(n137), .B(n473), .Q(n135) );
  INV2 U533 ( .A(n137), .Q(n471) );
  INV1 U534 ( .A(n176), .Q(n491) );
  XNR22 U535 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U536 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND22 U537 ( .A(n111), .B(n55), .Q(n53) );
  XNR22 U538 ( .A(n24), .B(n196), .Q(SUM[14]) );
  INV2 U539 ( .A(n111), .Q(n468) );
  NAND22 U540 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND22 U541 ( .A(n509), .B(n256), .Q(n32) );
  OAI211 U542 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  NAND24 U543 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR21 U544 ( .A(n194), .B(n497), .Q(n190) );
  INV1 U545 ( .A(n194), .Q(n507) );
  NAND21 U546 ( .A(n514), .B(n245), .Q(n30) );
  NOR22 U547 ( .A(n241), .B(n244), .Q(n239) );
  INV1 U548 ( .A(n255), .Q(n509) );
  INV2 U549 ( .A(n266), .Q(n504) );
  NAND21 U550 ( .A(n501), .B(n266), .Q(n34) );
  NOR22 U551 ( .A(A[12]), .B(B[12]), .Q(n212) );
  NAND21 U552 ( .A(A[13]), .B(B[13]), .Q(n206) );
  INV3 U553 ( .A(n219), .Q(n486) );
  NAND20 U554 ( .A(n485), .B(n224), .Q(n27) );
  OAI211 U555 ( .A(n88), .B(n465), .C(n89), .Q(n85) );
  NOR22 U556 ( .A(n99), .B(n106), .Q(n97) );
  CLKIN0 U557 ( .A(n239), .Q(n515) );
  INV0 U558 ( .A(n244), .Q(n514) );
  AOI210 U559 ( .A(n478), .B(n135), .C(n136), .Q(n130) );
  INV0 U560 ( .A(n136), .Q(n470) );
  NAND21 U561 ( .A(n490), .B(n89), .Q(n12) );
  NAND22 U562 ( .A(n486), .B(n203), .Q(n197) );
  NAND20 U563 ( .A(n507), .B(n195), .Q(n24) );
  INV0 U564 ( .A(n171), .Q(n492) );
  XOR21 U565 ( .A(n30), .B(n502), .Q(SUM[8]) );
  NAND22 U566 ( .A(n111), .B(n97), .Q(n91) );
  INV3 U567 ( .A(n5), .Q(n460) );
  NAND20 U568 ( .A(n239), .B(n488), .Q(n226) );
  INV0 U569 ( .A(n185), .Q(n494) );
  NAND20 U570 ( .A(n171), .B(n482), .Q(n158) );
  CLKIN0 U571 ( .A(n173), .Q(n495) );
  NAND20 U572 ( .A(n242), .B(n516), .Q(n29) );
  CLKIN0 U573 ( .A(n205), .Q(n496) );
  INV0 U574 ( .A(n117), .Q(n467) );
  NAND20 U575 ( .A(n467), .B(n118), .Q(n15) );
  INV0 U576 ( .A(n231), .Q(n487) );
  INV0 U577 ( .A(n155), .Q(n479) );
  CLKIN0 U578 ( .A(n252), .Q(n508) );
  INV0 U579 ( .A(n265), .Q(n501) );
  NAND20 U580 ( .A(A[20]), .B(B[20]), .Q(n432) );
  NAND20 U581 ( .A(A[20]), .B(B[20]), .Q(n431) );
  NAND20 U582 ( .A(n423), .B(n431), .Q(n18) );
  NOR20 U583 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR20 U584 ( .A(n46), .B(n6), .Q(n44) );
  INV0 U585 ( .A(n99), .Q(n511) );
  NOR21 U586 ( .A(n88), .B(n462), .Q(n84) );
  NAND20 U587 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U588 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U589 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U590 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV3 U591 ( .A(n19), .Q(n477) );
  NAND22 U592 ( .A(n480), .B(n135), .Q(n129) );
  NAND22 U593 ( .A(n480), .B(n122), .Q(n120) );
  INV0 U594 ( .A(n172), .Q(n493) );
  AOI210 U595 ( .A(n172), .B(n482), .C(n483), .Q(n159) );
  NAND22 U596 ( .A(n491), .B(n177), .Q(n22) );
  XOR21 U597 ( .A(n32), .B(n257), .Q(SUM[6]) );
  INV3 U598 ( .A(n126), .Q(n469) );
  NAND22 U599 ( .A(n496), .B(n206), .Q(n25) );
  NAND22 U600 ( .A(n494), .B(n186), .Q(n23) );
  NAND22 U601 ( .A(n471), .B(n138), .Q(n17) );
  NAND22 U602 ( .A(n508), .B(n253), .Q(n31) );
  NOR21 U603 ( .A(n126), .B(n472), .Q(n122) );
  NAND22 U604 ( .A(n479), .B(n156), .Q(n19) );
  NAND20 U605 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U606 ( .A(n212), .Q(n500) );
  INV3 U607 ( .A(n6), .Q(n459) );
  INV3 U608 ( .A(n60), .Q(n454) );
  XOR21 U609 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND22 U610 ( .A(n510), .B(n261), .Q(n33) );
  AOI211 U611 ( .A(n505), .B(n501), .C(n504), .Q(n262) );
  INV0 U612 ( .A(n260), .Q(n510) );
  NAND22 U613 ( .A(A[10]), .B(B[10]), .Q(n231) );
  INV3 U614 ( .A(n432), .Q(n475) );
  INV3 U615 ( .A(n12), .Q(n489) );
  NAND22 U616 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND22 U617 ( .A(A[9]), .B(B[9]), .Q(n242) );
  INV3 U618 ( .A(n59), .Q(n456) );
  INV3 U619 ( .A(n277), .Q(n519) );
  NAND22 U620 ( .A(n457), .B(n71), .Q(n10) );
  INV3 U621 ( .A(n70), .Q(n457) );
  NAND22 U622 ( .A(n455), .B(n62), .Q(n9) );
  INV3 U623 ( .A(n61), .Q(n455) );
  NAND22 U624 ( .A(n452), .B(n51), .Q(n8) );
  NAND20 U625 ( .A(n511), .B(n100), .Q(n13) );
  AOI210 U626 ( .A(n60), .B(n452), .C(n453), .Q(n47) );
  INV3 U627 ( .A(n51), .Q(n453) );
  NAND22 U628 ( .A(n458), .B(n80), .Q(n11) );
  NOR21 U629 ( .A(n61), .B(n70), .Q(n59) );
  INV3 U630 ( .A(n97), .Q(n462) );
  INV3 U631 ( .A(n88), .Q(n490) );
  NAND20 U632 ( .A(n59), .B(n452), .Q(n46) );
  XNR21 U633 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND20 U634 ( .A(n506), .B(n272), .Q(n35) );
  INV3 U635 ( .A(n271), .Q(n506) );
  XOR21 U636 ( .A(n36), .B(n519), .Q(SUM[2]) );
  NAND22 U637 ( .A(n512), .B(n275), .Q(n36) );
  INV3 U638 ( .A(n274), .Q(n512) );
  XOR21 U639 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U640 ( .A(n520), .B(n279), .Q(n37) );
  INV3 U641 ( .A(n278), .Q(n520) );
  XNR21 U642 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U643 ( .A(n451), .B(n40), .Q(n7) );
  NAND22 U644 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND21 U645 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NOR22 U646 ( .A(B[25]), .B(A[25]), .Q(n99) );
  INV3 U647 ( .A(n50), .Q(n452) );
  NOR20 U648 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NOR20 U649 ( .A(B[2]), .B(A[2]), .Q(n274) );
  INV3 U650 ( .A(n39), .Q(n451) );
  NOR21 U651 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND20 U652 ( .A(A[2]), .B(B[2]), .Q(n275) );
  INV3 U653 ( .A(n38), .Q(SUM[0]) );
  NAND22 U654 ( .A(n518), .B(n281), .Q(n38) );
  INV3 U655 ( .A(n280), .Q(n518) );
  NOR20 U656 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U657 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NOR20 U658 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND20 U659 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND22 U660 ( .A(n90), .B(n12), .Q(n426) );
  AOI210 U661 ( .A(n435), .B(n44), .C(n45), .Q(n43) );
  AOI210 U662 ( .A(n437), .B(n488), .C(n487), .Q(n227) );
  OAI210 U663 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  NOR21 U664 ( .A(B[24]), .B(A[24]), .Q(n106) );
endmodule


module adder_42 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1, n3, n4;

  adder_42_DW01_add_0 add_16 ( .A({A[31:21], n4, A[19:0]}), .B(B), .CI(n1), 
        .SUM(O) );
  INV4 U1 ( .A(A[20]), .Q(n3) );
  CLKIN6 U2 ( .A(n3), .Q(n4) );
  LOGIC0 U3 ( .Q(n1) );
endmodule


module adder_41_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n50,
         n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n418, n423, n426,
         n441, n512, n518, n519, n522, n526, n535, n602, n604, n618, n621,
         n698, n776, n785, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n936;

  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U490 ( .A(n241), .B(n245), .C(n242), .Q(n240) );
  AOI212 U522 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U540 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U544 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U357 ( .A(n176), .B(n863), .C(n177), .Q(n175) );
  OAI212 U462 ( .A(n5), .B(n892), .C(n894), .Q(n56) );
  NOR24 U466 ( .A(B[22]), .B(A[22]), .Q(n126) );
  OAI212 U474 ( .A(n113), .B(n860), .C(n114), .Q(n112) );
  OAI212 U509 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U567 ( .A(n152), .B(n113), .C(n114), .Q(n698) );
  NOR24 U427 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR24 U476 ( .A(A[17]), .B(B[17]), .Q(n173) );
  OAI212 U498 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  NOR24 U510 ( .A(B[25]), .B(A[25]), .Q(n99) );
  AOI212 U555 ( .A(n602), .B(n77), .C(n78), .Q(n604) );
  OAI212 U562 ( .A(n82), .B(n863), .C(n83), .Q(n81) );
  OAI212 U437 ( .A(n158), .B(n863), .C(n159), .Q(n157) );
  OAI212 U438 ( .A(n870), .B(n863), .C(n867), .Q(n164) );
  OAI210 U349 ( .A(n197), .B(n924), .C(n198), .Q(n196) );
  INV2 U350 ( .A(n145), .Q(n903) );
  NOR24 U351 ( .A(n117), .B(n126), .Q(n115) );
  NAND26 U352 ( .A(n618), .B(n80), .Q(n78) );
  INV6 U353 ( .A(n112), .Q(n865) );
  INV1 U354 ( .A(n136), .Q(n879) );
  NAND23 U355 ( .A(n441), .B(n65), .Q(n63) );
  NOR24 U356 ( .A(n223), .B(n230), .Q(n221) );
  NOR22 U358 ( .A(n260), .B(n265), .Q(n258) );
  CLKIN3 U359 ( .A(n860), .Q(n864) );
  AOI212 U360 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR22 U361 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR24 U362 ( .A(A[23]), .B(B[23]), .Q(n117) );
  NOR24 U363 ( .A(A[15]), .B(B[15]), .Q(n185) );
  NOR23 U364 ( .A(B[24]), .B(A[24]), .Q(n106) );
  OAI212 U365 ( .A(n126), .B(n879), .C(n127), .Q(n123) );
  XNR22 U366 ( .A(n90), .B(n862), .Q(SUM[26]) );
  NOR24 U367 ( .A(n865), .B(n887), .Q(n526) );
  XNR22 U368 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NOR24 U369 ( .A(A[18]), .B(B[18]), .Q(n162) );
  NOR23 U370 ( .A(n155), .B(n162), .Q(n153) );
  NAND26 U371 ( .A(n621), .B(n174), .Q(n172) );
  BUF12 U372 ( .A(n698), .Q(n859) );
  NAND23 U373 ( .A(n239), .B(n221), .Q(n219) );
  NAND26 U374 ( .A(n153), .B(n171), .Q(n151) );
  NAND21 U375 ( .A(n871), .B(n902), .Q(n140) );
  AOI211 U376 ( .A(n864), .B(n135), .C(n861), .Q(n130) );
  INV0 U377 ( .A(n244), .Q(n923) );
  NOR22 U378 ( .A(n241), .B(n244), .Q(n239) );
  OAI211 U379 ( .A(n140), .B(n863), .C(n141), .Q(n139) );
  NOR23 U380 ( .A(n194), .B(n185), .Q(n183) );
  NAND22 U381 ( .A(A[26]), .B(B[26]), .Q(n89) );
  INV3 U382 ( .A(n97), .Q(n885) );
  NAND22 U383 ( .A(n905), .B(n868), .Q(n518) );
  NAND23 U384 ( .A(n906), .B(n866), .Q(n621) );
  NAND22 U385 ( .A(n111), .B(n66), .Q(n64) );
  NOR22 U386 ( .A(n70), .B(n6), .Q(n66) );
  NOR23 U387 ( .A(A[27]), .B(B[27]), .Q(n79) );
  NOR23 U388 ( .A(A[21]), .B(B[21]), .Q(n137) );
  NOR23 U389 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NOR21 U390 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR22 U391 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR23 U392 ( .A(A[11]), .B(B[11]), .Q(n223) );
  NAND23 U393 ( .A(n512), .B(n206), .Q(n204) );
  NOR23 U394 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR22 U395 ( .A(n252), .B(n255), .Q(n250) );
  NAND22 U396 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NOR21 U397 ( .A(n126), .B(n881), .Q(n122) );
  NOR22 U398 ( .A(n88), .B(n885), .Q(n84) );
  NAND23 U399 ( .A(n776), .B(n74), .Q(n72) );
  NAND22 U400 ( .A(n876), .B(n907), .Q(n426) );
  NAND23 U401 ( .A(n54), .B(n535), .Q(n52) );
  NAND22 U402 ( .A(n891), .B(n62), .Q(n9) );
  NAND22 U403 ( .A(n519), .B(n518), .Q(SUM[17]) );
  XNR21 U404 ( .A(n16), .B(n128), .Q(SUM[22]) );
  AOI212 U405 ( .A(n172), .B(n153), .C(n154), .Q(n860) );
  CLKIN2 U406 ( .A(n203), .Q(n912) );
  INV3 U407 ( .A(n879), .Q(n861) );
  NAND21 U408 ( .A(n917), .B(n203), .Q(n197) );
  NAND24 U409 ( .A(n203), .B(n183), .Q(n181) );
  INV3 U410 ( .A(n247), .Q(n924) );
  NAND21 U411 ( .A(A[3]), .B(B[3]), .Q(n272) );
  OAI212 U412 ( .A(n120), .B(n863), .C(n121), .Q(n119) );
  INV0 U413 ( .A(n61), .Q(n891) );
  NAND22 U414 ( .A(B[9]), .B(A[9]), .Q(n242) );
  OAI212 U415 ( .A(n241), .B(n245), .C(n242), .Q(n785) );
  NAND24 U416 ( .A(n522), .B(n47), .Q(n45) );
  NAND21 U417 ( .A(B[21]), .B(A[21]), .Q(n138) );
  NOR22 U418 ( .A(n173), .B(n176), .Q(n171) );
  NOR24 U419 ( .A(n181), .B(n219), .Q(n179) );
  NAND24 U420 ( .A(n897), .B(n898), .Q(n618) );
  NAND21 U421 ( .A(B[23]), .B(A[23]), .Q(n118) );
  OAI212 U422 ( .A(n129), .B(n863), .C(n130), .Q(n128) );
  CLKIN6 U423 ( .A(n173), .Q(n906) );
  AOI211 U424 ( .A(n60), .B(n895), .C(n896), .Q(n47) );
  NAND21 U425 ( .A(n895), .B(n51), .Q(n8) );
  NAND21 U426 ( .A(A[30]), .B(B[30]), .Q(n51) );
  AOI211 U428 ( .A(n864), .B(n902), .C(n903), .Q(n141) );
  INV3 U429 ( .A(n135), .Q(n881) );
  NAND26 U430 ( .A(n135), .B(n115), .Q(n113) );
  NOR23 U431 ( .A(n144), .B(n137), .Q(n135) );
  INV4 U432 ( .A(n604), .Q(n889) );
  NAND24 U433 ( .A(n893), .B(n889), .Q(n522) );
  INV12 U434 ( .A(n863), .Q(n907) );
  NAND24 U435 ( .A(n59), .B(n895), .Q(n46) );
  INV6 U436 ( .A(n50), .Q(n895) );
  AOI212 U439 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND21 U440 ( .A(n871), .B(n135), .Q(n129) );
  OAI212 U441 ( .A(n604), .B(n70), .C(n71), .Q(n67) );
  NAND22 U442 ( .A(A[17]), .B(B[17]), .Q(n174) );
  AOI211 U443 ( .A(n859), .B(n886), .C(n889), .Q(n74) );
  OAI211 U444 ( .A(n107), .B(n99), .C(n100), .Q(n602) );
  NAND22 U445 ( .A(B[25]), .B(A[25]), .Q(n100) );
  NOR24 U446 ( .A(B[26]), .B(A[26]), .Q(n88) );
  OAI212 U447 ( .A(n88), .B(n890), .C(n89), .Q(n85) );
  INV2 U448 ( .A(n51), .Q(n896) );
  NAND22 U449 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NOR24 U450 ( .A(n892), .B(n6), .Q(n55) );
  OAI212 U451 ( .A(n91), .B(n863), .C(n92), .Q(n90) );
  NAND20 U452 ( .A(n902), .B(n145), .Q(n18) );
  INV1 U453 ( .A(n144), .Q(n902) );
  NAND22 U454 ( .A(n111), .B(n97), .Q(n91) );
  NAND22 U455 ( .A(n111), .B(n44), .Q(n42) );
  NAND24 U456 ( .A(n907), .B(n874), .Q(n535) );
  NAND21 U457 ( .A(n111), .B(n84), .Q(n82) );
  NAND21 U458 ( .A(n111), .B(n886), .Q(n73) );
  INV2 U459 ( .A(n220), .Q(n915) );
  NAND24 U460 ( .A(n426), .B(n43), .Q(n41) );
  NOR24 U461 ( .A(n45), .B(n526), .Q(n43) );
  AOI212 U463 ( .A(n859), .B(n84), .C(n85), .Q(n83) );
  OAI212 U464 ( .A(n863), .B(n102), .C(n103), .Q(n101) );
  NAND21 U465 ( .A(n111), .B(n884), .Q(n102) );
  XNR22 U467 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR22 U468 ( .A(n9), .B(n63), .Q(SUM[29]) );
  AOI211 U469 ( .A(n112), .B(n97), .C(n98), .Q(n92) );
  XNR22 U470 ( .A(n7), .B(n41), .Q(SUM[31]) );
  XNR22 U471 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NOR24 U472 ( .A(n61), .B(n70), .Q(n59) );
  INV0 U473 ( .A(n70), .Q(n899) );
  NOR24 U475 ( .A(B[28]), .B(A[28]), .Q(n70) );
  INV3 U477 ( .A(n44), .Q(n887) );
  NOR23 U478 ( .A(n46), .B(n6), .Q(n44) );
  NOR22 U479 ( .A(B[30]), .B(A[30]), .Q(n50) );
  OAI210 U480 ( .A(n173), .B(n177), .C(n174), .Q(n423) );
  NOR22 U481 ( .A(n271), .B(n274), .Q(n269) );
  OAI210 U482 ( .A(n274), .B(n933), .C(n275), .Q(n273) );
  OAI211 U483 ( .A(n872), .B(n863), .C(n865), .Q(n108) );
  INV1 U484 ( .A(n111), .Q(n872) );
  OAI211 U485 ( .A(n194), .B(n910), .C(n195), .Q(n191) );
  NAND22 U486 ( .A(A[14]), .B(B[14]), .Q(n195) );
  OAI211 U487 ( .A(n208), .B(n924), .C(n209), .Q(n207) );
  INV0 U488 ( .A(n155), .Q(n904) );
  NOR24 U489 ( .A(A[19]), .B(B[19]), .Q(n155) );
  OAI212 U491 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND21 U492 ( .A(A[29]), .B(B[29]), .Q(n62) );
  CLKIN2 U493 ( .A(n60), .Q(n894) );
  XOR20 U494 ( .A(n30), .B(n924), .Q(SUM[8]) );
  OAI210 U495 ( .A(n219), .B(n924), .C(n220), .Q(n214) );
  OAI210 U496 ( .A(n244), .B(n924), .C(n245), .Q(n243) );
  OAI210 U497 ( .A(n226), .B(n924), .C(n227), .Q(n225) );
  OAI210 U499 ( .A(n922), .B(n924), .C(n920), .Q(n232) );
  OAI211 U500 ( .A(n924), .B(n188), .C(n189), .Q(n187) );
  NAND22 U501 ( .A(A[20]), .B(B[20]), .Q(n145) );
  INV1 U502 ( .A(n46), .Q(n893) );
  AOI211 U503 ( .A(n859), .B(n55), .C(n56), .Q(n54) );
  AOI212 U504 ( .A(n859), .B(n884), .C(n888), .Q(n103) );
  NOR24 U505 ( .A(n88), .B(n79), .Q(n77) );
  CLKIN6 U506 ( .A(n79), .Q(n898) );
  INV6 U507 ( .A(n6), .Q(n886) );
  NAND28 U508 ( .A(n77), .B(n97), .Q(n6) );
  NOR24 U511 ( .A(B[29]), .B(A[29]), .Q(n61) );
  AOI211 U512 ( .A(n864), .B(n122), .C(n123), .Q(n121) );
  NAND22 U513 ( .A(B[13]), .B(A[13]), .Q(n206) );
  AOI211 U514 ( .A(n859), .B(n66), .C(n67), .Q(n65) );
  NAND24 U515 ( .A(B[18]), .B(A[18]), .Q(n163) );
  INV2 U516 ( .A(n163), .Q(n877) );
  AOI211 U517 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U518 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  NAND21 U519 ( .A(B[19]), .B(A[19]), .Q(n156) );
  NAND24 U520 ( .A(B[22]), .B(A[22]), .Q(n127) );
  NAND21 U521 ( .A(B[15]), .B(A[15]), .Q(n186) );
  OAI212 U523 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U524 ( .A(n137), .B(n145), .C(n138), .Q(n136) );
  NOR24 U525 ( .A(n99), .B(n106), .Q(n97) );
  NOR24 U526 ( .A(n113), .B(n151), .Q(n111) );
  OAI211 U527 ( .A(n151), .B(n863), .C(n860), .Q(n146) );
  AOI212 U528 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  NAND22 U529 ( .A(n899), .B(n71), .Q(n10) );
  NAND22 U530 ( .A(A[27]), .B(B[27]), .Q(n80) );
  OAI211 U531 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI211 U532 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NAND22 U533 ( .A(n926), .B(n256), .Q(n32) );
  NAND21 U534 ( .A(A[6]), .B(B[6]), .Q(n256) );
  INV0 U535 ( .A(n171), .Q(n870) );
  NAND22 U536 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NOR22 U537 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR24 U538 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND22 U539 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NOR22 U541 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR22 U542 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND22 U543 ( .A(n917), .B(n190), .Q(n188) );
  INV1 U545 ( .A(n98), .Q(n890) );
  INV3 U546 ( .A(n59), .Q(n892) );
  AOI211 U547 ( .A(n915), .B(n190), .C(n191), .Q(n189) );
  AOI210 U548 ( .A(n785), .B(n919), .C(n918), .Q(n227) );
  NOR22 U549 ( .A(n205), .B(n212), .Q(n203) );
  CLKIN0 U550 ( .A(n423), .Q(n867) );
  CLKIN3 U551 ( .A(n205), .Q(n911) );
  CLKIN0 U552 ( .A(n204), .Q(n910) );
  NAND22 U553 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND21 U554 ( .A(B[11]), .B(A[11]), .Q(n224) );
  NAND26 U556 ( .A(B[16]), .B(A[16]), .Q(n177) );
  NAND22 U557 ( .A(B[12]), .B(A[12]), .Q(n213) );
  NAND22 U558 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U559 ( .A(n875), .B(n907), .Q(n441) );
  INV2 U560 ( .A(n64), .Q(n875) );
  AOI210 U561 ( .A(n915), .B(n203), .C(n204), .Q(n198) );
  AOI210 U563 ( .A(n915), .B(n914), .C(n913), .Q(n209) );
  NAND22 U564 ( .A(n917), .B(n914), .Q(n208) );
  CLKIN6 U565 ( .A(n175), .Q(n868) );
  AOI212 U566 ( .A(n115), .B(n136), .C(n116), .Q(n114) );
  NAND21 U568 ( .A(n871), .B(n122), .Q(n120) );
  AOI212 U569 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  AOI210 U570 ( .A(n930), .B(n929), .C(n928), .Q(n262) );
  INV0 U571 ( .A(n231), .Q(n918) );
  INV0 U572 ( .A(n212), .Q(n914) );
  INV0 U573 ( .A(n265), .Q(n929) );
  INV0 U574 ( .A(n274), .Q(n932) );
  INV0 U575 ( .A(n277), .Q(n933) );
  INV0 U576 ( .A(n278), .Q(n934) );
  NAND21 U577 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND21 U578 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND21 U579 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U580 ( .A(n39), .Q(n900) );
  NAND20 U581 ( .A(n932), .B(n275), .Q(n36) );
  XNR20 U582 ( .A(n34), .B(n930), .Q(SUM[4]) );
  NAND20 U583 ( .A(n934), .B(n279), .Q(n37) );
  INV3 U584 ( .A(n53), .Q(n874) );
  NAND22 U585 ( .A(n111), .B(n55), .Q(n53) );
  NAND22 U586 ( .A(n873), .B(n907), .Q(n776) );
  INV3 U587 ( .A(n73), .Q(n873) );
  INV3 U588 ( .A(n42), .Q(n876) );
  INV3 U589 ( .A(n219), .Q(n917) );
  INV3 U590 ( .A(n151), .Q(n871) );
  NAND22 U591 ( .A(n21), .B(n175), .Q(n519) );
  INV3 U592 ( .A(n239), .Q(n922) );
  INV3 U593 ( .A(n785), .Q(n920) );
  AOI210 U594 ( .A(n930), .B(n258), .C(n259), .Q(n418) );
  INV3 U595 ( .A(n268), .Q(n930) );
  INV3 U596 ( .A(n21), .Q(n905) );
  NAND20 U597 ( .A(n171), .B(n878), .Q(n158) );
  AOI210 U598 ( .A(n423), .B(n878), .C(n877), .Q(n159) );
  INV3 U599 ( .A(n107), .Q(n888) );
  INV3 U600 ( .A(n89), .Q(n897) );
  NAND22 U601 ( .A(n258), .B(n250), .Q(n248) );
  AOI210 U602 ( .A(n930), .B(n258), .C(n259), .Q(n257) );
  NAND20 U603 ( .A(n239), .B(n919), .Q(n226) );
  NOR21 U604 ( .A(n194), .B(n912), .Q(n190) );
  INV3 U605 ( .A(n266), .Q(n928) );
  NAND22 U606 ( .A(n913), .B(n911), .Q(n512) );
  NAND20 U607 ( .A(n906), .B(n174), .Q(n21) );
  INV3 U608 ( .A(n106), .Q(n884) );
  INV3 U609 ( .A(n162), .Q(n878) );
  INV0 U610 ( .A(n194), .Q(n909) );
  INV0 U611 ( .A(n126), .Q(n882) );
  INV0 U612 ( .A(n241), .Q(n921) );
  INV0 U613 ( .A(n99), .Q(n901) );
  INV3 U614 ( .A(n177), .Q(n866) );
  INV3 U615 ( .A(n260), .Q(n927) );
  INV3 U616 ( .A(n255), .Q(n926) );
  INV3 U617 ( .A(n213), .Q(n913) );
  INV0 U618 ( .A(n117), .Q(n883) );
  INV3 U619 ( .A(n252), .Q(n925) );
  INV0 U620 ( .A(n185), .Q(n908) );
  INV0 U621 ( .A(n223), .Q(n916) );
  INV0 U622 ( .A(n176), .Q(n869) );
  INV3 U623 ( .A(n137), .Q(n880) );
  NAND22 U624 ( .A(n931), .B(n272), .Q(n35) );
  INV3 U625 ( .A(n271), .Q(n931) );
  NOR23 U626 ( .A(A[12]), .B(B[12]), .Q(n212) );
  NOR21 U627 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR23 U628 ( .A(A[13]), .B(B[13]), .Q(n205) );
  NOR21 U629 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U630 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U631 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND22 U632 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NOR21 U633 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U634 ( .A(n280), .Q(n936) );
  NOR21 U635 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U636 ( .A(n900), .B(n40), .Q(n7) );
  XNR21 U637 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NAND20 U638 ( .A(n901), .B(n100), .Q(n13) );
  XNR20 U639 ( .A(B[26]), .B(A[26]), .Q(n862) );
  XNR21 U640 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U641 ( .A(n156), .B(n904), .Q(n19) );
  XNR21 U642 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND20 U643 ( .A(n882), .B(n127), .Q(n16) );
  XNR21 U644 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND20 U645 ( .A(n883), .B(n118), .Q(n15) );
  NAND20 U646 ( .A(n898), .B(n80), .Q(n11) );
  XNR21 U647 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND20 U648 ( .A(n884), .B(n107), .Q(n14) );
  XNR21 U649 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND20 U650 ( .A(n878), .B(n163), .Q(n20) );
  XNR21 U651 ( .A(n17), .B(n139), .Q(SUM[21]) );
  NAND20 U652 ( .A(n880), .B(n138), .Q(n17) );
  XOR20 U653 ( .A(n22), .B(n863), .Q(SUM[16]) );
  NAND20 U654 ( .A(n869), .B(n177), .Q(n22) );
  XNR21 U655 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U656 ( .A(n909), .B(n195), .Q(n24) );
  XNR21 U657 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U658 ( .A(n911), .B(n206), .Q(n25) );
  XNR21 U659 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U660 ( .A(n916), .B(n224), .Q(n27) );
  XNR21 U661 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U662 ( .A(n919), .B(n231), .Q(n28) );
  NAND20 U663 ( .A(n923), .B(n245), .Q(n30) );
  NAND20 U664 ( .A(n929), .B(n266), .Q(n34) );
  XOR21 U665 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND20 U666 ( .A(n927), .B(n261), .Q(n33) );
  XNR21 U667 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U668 ( .A(n908), .B(n186), .Q(n23) );
  XNR21 U669 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U670 ( .A(n213), .B(n914), .Q(n26) );
  XNR21 U671 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U672 ( .A(n921), .B(n242), .Q(n29) );
  XOR21 U673 ( .A(n32), .B(n418), .Q(SUM[6]) );
  XNR21 U674 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U675 ( .A(n925), .B(n253), .Q(n31) );
  XOR21 U676 ( .A(n281), .B(n37), .Q(SUM[1]) );
  XNR21 U677 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XOR21 U678 ( .A(n36), .B(n933), .Q(SUM[2]) );
  INV3 U679 ( .A(n38), .Q(SUM[0]) );
  NAND22 U680 ( .A(n936), .B(n281), .Q(n38) );
  CLKIN3 U681 ( .A(n230), .Q(n919) );
  BUF15 U682 ( .A(n178), .Q(n863) );
endmodule


module adder_41 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_41_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module reg_13 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30,
         n32, n35, n47, n49, n51, n53, n55, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n58, n59, n60, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n107, n108, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393;

  DF3 Dout_reg_16_ ( .D(n76), .C(Clk), .Q(Dout[16]), .QN(n14) );
  DF3 Dout_reg_15_ ( .D(n77), .C(Clk), .Q(Dout[15]), .QN(n12) );
  DF3 Dout_reg_14_ ( .D(n78), .C(Clk), .Q(Dout[14]), .QN(n10) );
  DF3 Dout_reg_13_ ( .D(n79), .C(Clk), .Q(Dout[13]), .QN(n8) );
  DF3 Dout_reg_12_ ( .D(n80), .C(Clk), .Q(Dout[12]), .QN(n6) );
  DF3 Dout_reg_11_ ( .D(n81), .C(Clk), .Q(Dout[11]), .QN(n4) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n58) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n59) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n85) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n84) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n83) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n82) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n88) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n87) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n89) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n60) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n86) );
  OAI222 U3 ( .A(n86), .B(n358), .C(n360), .D(n392), .Q(n99) );
  OAI222 U4 ( .A(n87), .B(n358), .C(n359), .D(n390), .Q(n98) );
  OAI222 U5 ( .A(n88), .B(n358), .C(n107), .D(n391), .Q(n97) );
  OAI222 U6 ( .A(n82), .B(n358), .C(n360), .D(n389), .Q(n96) );
  OAI222 U7 ( .A(n83), .B(n358), .C(n359), .D(n388), .Q(n95) );
  OAI222 U8 ( .A(n84), .B(n358), .C(n107), .D(n387), .Q(n94) );
  OAI222 U9 ( .A(n85), .B(n358), .C(n360), .D(n386), .Q(n93) );
  OAI222 U10 ( .A(n59), .B(n358), .C(n359), .D(n385), .Q(n92) );
  OAI222 U11 ( .A(n60), .B(n358), .C(n107), .D(n384), .Q(n91) );
  OAI222 U12 ( .A(n58), .B(n358), .C(n360), .D(n383), .Q(n90) );
  OAI222 U13 ( .A(n4), .B(n358), .C(n359), .D(n382), .Q(n81) );
  OAI222 U14 ( .A(n6), .B(n358), .C(n107), .D(n381), .Q(n80) );
  OAI222 U15 ( .A(n8), .B(n358), .C(n360), .D(n380), .Q(n79) );
  OAI222 U16 ( .A(n10), .B(n358), .C(n359), .D(n379), .Q(n78) );
  OAI222 U17 ( .A(n12), .B(n358), .C(n107), .D(n378), .Q(n77) );
  OAI222 U18 ( .A(n14), .B(n358), .C(n360), .D(n363), .Q(n76) );
  OAI222 U19 ( .A(n16), .B(n358), .C(n359), .D(n362), .Q(n75) );
  OAI222 U20 ( .A(n18), .B(n358), .C(n107), .D(n364), .Q(n74) );
  OAI222 U21 ( .A(n20), .B(n358), .C(n360), .D(n365), .Q(n73) );
  OAI222 U22 ( .A(n22), .B(n358), .C(n359), .D(n377), .Q(n72) );
  OAI222 U23 ( .A(n24), .B(n358), .C(n107), .D(n374), .Q(n71) );
  OAI222 U24 ( .A(n26), .B(n358), .C(n360), .D(n373), .Q(n70) );
  OAI222 U25 ( .A(n28), .B(n358), .C(n359), .D(n375), .Q(n69) );
  OAI222 U26 ( .A(n30), .B(n358), .C(n107), .D(n376), .Q(n68) );
  OAI222 U27 ( .A(n32), .B(n358), .C(n360), .D(n367), .Q(n67) );
  OAI222 U28 ( .A(n35), .B(n358), .C(n359), .D(n372), .Q(n66) );
  OAI222 U29 ( .A(n47), .B(n358), .C(n107), .D(n366), .Q(n65) );
  OAI222 U30 ( .A(n49), .B(n358), .C(n360), .D(n368), .Q(n64) );
  OAI222 U31 ( .A(n51), .B(n358), .C(n359), .D(n370), .Q(n63) );
  OAI222 U32 ( .A(n53), .B(n358), .C(n107), .D(n369), .Q(n62) );
  OAI222 U33 ( .A(n55), .B(n358), .C(n360), .D(n371), .Q(n61) );
  OAI222 U34 ( .A(n89), .B(n358), .C(n359), .D(n393), .Q(n100) );
  DF1 Dout_reg_21_ ( .D(n71), .C(Clk), .Q(Dout[21]), .QN(n24) );
  DF1 Dout_reg_18_ ( .D(n74), .C(Clk), .Q(Dout[18]), .QN(n18) );
  DF1 Dout_reg_20_ ( .D(n72), .C(Clk), .Q(Dout[20]), .QN(n22) );
  DF1 Dout_reg_17_ ( .D(n75), .C(Clk), .Q(Dout[17]), .QN(n16) );
  DF1 Dout_reg_31_ ( .D(n61), .C(Clk), .Q(Dout[31]), .QN(n55) );
  DF1 Dout_reg_23_ ( .D(n69), .C(Clk), .Q(Dout[23]), .QN(n28) );
  DF1 Dout_reg_22_ ( .D(n70), .C(Clk), .Q(Dout[22]), .QN(n26) );
  DF1 Dout_reg_19_ ( .D(n73), .C(Clk), .Q(Dout[19]), .QN(n20) );
  DF1 Dout_reg_24_ ( .D(n68), .C(Clk), .Q(Dout[24]), .QN(n30) );
  DF1 Dout_reg_28_ ( .D(n64), .C(Clk), .Q(Dout[28]), .QN(n49) );
  DF1 Dout_reg_27_ ( .D(n65), .C(Clk), .Q(Dout[27]), .QN(n47) );
  DF1 Dout_reg_26_ ( .D(n66), .C(Clk), .Q(Dout[26]), .QN(n35) );
  DF1 Dout_reg_30_ ( .D(n62), .C(Clk), .Q(Dout[30]), .QN(n53) );
  DF1 Dout_reg_29_ ( .D(n63), .C(Clk), .Q(Dout[29]), .QN(n51) );
  DF1 Dout_reg_25_ ( .D(n67), .C(Clk), .Q(Dout[25]), .QN(n32) );
  INV4 U35 ( .A(Din[29]), .Q(n370) );
  INV4 U36 ( .A(Din[26]), .Q(n372) );
  INV3 U37 ( .A(Din[28]), .Q(n368) );
  INV4 U38 ( .A(Din[27]), .Q(n366) );
  INV4 U39 ( .A(Din[30]), .Q(n369) );
  INV3 U40 ( .A(Din[31]), .Q(n371) );
  INV2 U41 ( .A(Din[16]), .Q(n363) );
  INV2 U42 ( .A(Din[12]), .Q(n381) );
  CLKIN3 U43 ( .A(Din[8]), .Q(n385) );
  INV2 U44 ( .A(Din[24]), .Q(n376) );
  INV2 U45 ( .A(Din[19]), .Q(n365) );
  INV2 U46 ( .A(Din[23]), .Q(n375) );
  INV2 U47 ( .A(Din[22]), .Q(n373) );
  INV2 U48 ( .A(Din[20]), .Q(n377) );
  INV3 U49 ( .A(Din[17]), .Q(n362) );
  INV2 U50 ( .A(Din[14]), .Q(n379) );
  INV2 U51 ( .A(Din[13]), .Q(n380) );
  INV2 U52 ( .A(Din[10]), .Q(n383) );
  INV2 U53 ( .A(Din[11]), .Q(n382) );
  INV2 U54 ( .A(Din[7]), .Q(n386) );
  INV2 U55 ( .A(Din[21]), .Q(n374) );
  INV2 U56 ( .A(Din[18]), .Q(n364) );
  INV2 U57 ( .A(Din[15]), .Q(n378) );
  INV2 U58 ( .A(Din[9]), .Q(n384) );
  CLKIN3 U59 ( .A(Din[6]), .Q(n387) );
  NAND22 U60 ( .A(n361), .B(n358), .Q(n359) );
  NAND22 U61 ( .A(n361), .B(n358), .Q(n360) );
  NAND22 U62 ( .A(n361), .B(n358), .Q(n107) );
  INV3 U63 ( .A(Reset), .Q(n361) );
  INV3 U64 ( .A(n108), .Q(n358) );
  INV3 U65 ( .A(Din[25]), .Q(n367) );
  INV3 U66 ( .A(Din[4]), .Q(n389) );
  INV3 U67 ( .A(Din[5]), .Q(n388) );
  INV3 U68 ( .A(Din[3]), .Q(n391) );
  INV3 U69 ( .A(Din[1]), .Q(n392) );
  INV3 U70 ( .A(Din[2]), .Q(n390) );
  INV3 U71 ( .A(Din[0]), .Q(n393) );
  NOR20 U72 ( .A(Load), .B(Reset), .Q(n108) );
endmodule


module reg_12 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32,
         n35, n47, n49, n51, n53, n55, n57, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n58, n59, n60, n61, n62, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n105, n106, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395;

  DF3 Dout_reg_16_ ( .D(n78), .C(Clk), .Q(Dout[16]), .QN(n16) );
  DF3 Dout_reg_15_ ( .D(n79), .C(Clk), .Q(Dout[15]), .QN(n14) );
  DF3 Dout_reg_14_ ( .D(n80), .C(Clk), .Q(Dout[14]), .QN(n12) );
  DF3 Dout_reg_12_ ( .D(n82), .C(Clk), .Q(Dout[12]), .QN(n8) );
  DF3 Dout_reg_11_ ( .D(n83), .C(Clk), .Q(Dout[11]), .QN(n6) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n58) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n59) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n85) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n84) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n62) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n61) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n87) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n89) );
  DF3 Dout_reg_13_ ( .D(n81), .C(Clk), .Q(Dout[13]), .QN(n10) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n60) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n88) );
  DF3 Dout_reg_26_ ( .D(n68), .C(Clk), .Q(Dout[26]), .QN(n47) );
  OAI222 U3 ( .A(n86), .B(n360), .C(n362), .D(n394), .Q(n99) );
  OAI222 U4 ( .A(n87), .B(n360), .C(n361), .D(n392), .Q(n98) );
  OAI222 U5 ( .A(n88), .B(n360), .C(n105), .D(n393), .Q(n97) );
  OAI222 U6 ( .A(n61), .B(n360), .C(n362), .D(n391), .Q(n96) );
  OAI222 U7 ( .A(n62), .B(n360), .C(n361), .D(n390), .Q(n95) );
  OAI222 U8 ( .A(n84), .B(n360), .C(n105), .D(n389), .Q(n94) );
  OAI222 U9 ( .A(n85), .B(n360), .C(n362), .D(n388), .Q(n93) );
  OAI222 U10 ( .A(n59), .B(n360), .C(n361), .D(n386), .Q(n92) );
  OAI222 U11 ( .A(n60), .B(n360), .C(n105), .D(n387), .Q(n91) );
  OAI222 U12 ( .A(n58), .B(n360), .C(n362), .D(n385), .Q(n90) );
  OAI222 U13 ( .A(n6), .B(n360), .C(n361), .D(n384), .Q(n83) );
  OAI222 U14 ( .A(n8), .B(n360), .C(n105), .D(n382), .Q(n82) );
  OAI222 U15 ( .A(n10), .B(n360), .C(n362), .D(n383), .Q(n81) );
  OAI222 U16 ( .A(n12), .B(n360), .C(n361), .D(n381), .Q(n80) );
  OAI222 U17 ( .A(n14), .B(n360), .C(n105), .D(n380), .Q(n79) );
  OAI222 U18 ( .A(n16), .B(n360), .C(n362), .D(n364), .Q(n78) );
  OAI222 U19 ( .A(n18), .B(n360), .C(n361), .D(n379), .Q(n77) );
  OAI222 U20 ( .A(n20), .B(n360), .C(n105), .D(n365), .Q(n76) );
  OAI222 U21 ( .A(n22), .B(n360), .C(n362), .D(n378), .Q(n75) );
  OAI222 U22 ( .A(n24), .B(n360), .C(n361), .D(n377), .Q(n74) );
  OAI222 U23 ( .A(n26), .B(n360), .C(n367), .D(n105), .Q(n73) );
  OAI222 U24 ( .A(n28), .B(n360), .C(n362), .D(n368), .Q(n72) );
  OAI222 U25 ( .A(n30), .B(n360), .C(n361), .D(n366), .Q(n71) );
  OAI222 U26 ( .A(n32), .B(n360), .C(n105), .D(n369), .Q(n70) );
  OAI222 U27 ( .A(n35), .B(n360), .C(n362), .D(n370), .Q(n69) );
  OAI222 U28 ( .A(n47), .B(n360), .C(n361), .D(n373), .Q(n68) );
  OAI222 U29 ( .A(n49), .B(n360), .C(n105), .D(n372), .Q(n67) );
  OAI222 U30 ( .A(n51), .B(n360), .C(n362), .D(n371), .Q(n66) );
  OAI222 U31 ( .A(n53), .B(n360), .C(n375), .D(n361), .Q(n65) );
  OAI222 U32 ( .A(n55), .B(n360), .C(n105), .D(n374), .Q(n64) );
  OAI222 U33 ( .A(n57), .B(n360), .C(n362), .D(n376), .Q(n63) );
  OAI222 U34 ( .A(n89), .B(n360), .C(n361), .D(n395), .Q(n100) );
  DF1 Dout_reg_27_ ( .D(n67), .C(Clk), .Q(Dout[27]), .QN(n49) );
  DF1 Dout_reg_23_ ( .D(n71), .C(Clk), .Q(Dout[23]), .QN(n30) );
  DF1 Dout_reg_22_ ( .D(n72), .C(Clk), .Q(Dout[22]), .QN(n28) );
  DF1 Dout_reg_20_ ( .D(n74), .C(Clk), .Q(Dout[20]), .QN(n24) );
  DF1 Dout_reg_18_ ( .D(n76), .C(Clk), .Q(Dout[18]), .QN(n20) );
  DF1 Dout_reg_31_ ( .D(n63), .C(Clk), .Q(Dout[31]), .QN(n57) );
  DF1 Dout_reg_30_ ( .D(n64), .C(Clk), .Q(Dout[30]), .QN(n55) );
  DF3 Dout_reg_29_ ( .D(n65), .C(Clk), .Q(Dout[29]), .QN(n53) );
  DF3 Dout_reg_28_ ( .D(n66), .C(Clk), .Q(Dout[28]), .QN(n51) );
  DF3 Dout_reg_24_ ( .D(n70), .C(Clk), .Q(Dout[24]), .QN(n32) );
  DF3 Dout_reg_25_ ( .D(n69), .C(Clk), .Q(Dout[25]), .QN(n35) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n86) );
  DF3 Dout_reg_21_ ( .D(n73), .C(Clk), .Q(Dout[21]), .QN(n26) );
  DF3 Dout_reg_17_ ( .D(n77), .C(Clk), .Q(Dout[17]), .QN(n18) );
  DF1 Dout_reg_19_ ( .D(n75), .C(Clk), .Q(Dout[19]), .QN(n22) );
  INV4 U35 ( .A(Din[31]), .Q(n376) );
  INV4 U36 ( .A(Din[30]), .Q(n374) );
  INV4 U37 ( .A(Din[25]), .Q(n370) );
  INV3 U38 ( .A(Din[21]), .Q(n367) );
  INV3 U39 ( .A(Din[29]), .Q(n375) );
  INV2 U40 ( .A(Din[7]), .Q(n388) );
  INV2 U41 ( .A(Din[4]), .Q(n391) );
  CLKIN3 U42 ( .A(Din[6]), .Q(n389) );
  INV3 U43 ( .A(Din[8]), .Q(n386) );
  INV2 U44 ( .A(Din[28]), .Q(n371) );
  INV2 U45 ( .A(Din[26]), .Q(n373) );
  INV2 U46 ( .A(Din[17]), .Q(n379) );
  INV2 U47 ( .A(Din[23]), .Q(n366) );
  INV2 U48 ( .A(Din[19]), .Q(n378) );
  INV2 U49 ( .A(Din[20]), .Q(n377) );
  INV2 U50 ( .A(Din[22]), .Q(n368) );
  INV2 U51 ( .A(Din[16]), .Q(n364) );
  INV2 U52 ( .A(Din[13]), .Q(n383) );
  INV2 U53 ( .A(Din[14]), .Q(n381) );
  INV2 U54 ( .A(Din[11]), .Q(n384) );
  INV2 U55 ( .A(Din[10]), .Q(n385) );
  INV2 U56 ( .A(Din[24]), .Q(n369) );
  INV2 U57 ( .A(Din[27]), .Q(n372) );
  INV2 U58 ( .A(Din[18]), .Q(n365) );
  INV2 U59 ( .A(Din[15]), .Q(n380) );
  INV2 U60 ( .A(Din[9]), .Q(n387) );
  INV2 U61 ( .A(Din[12]), .Q(n382) );
  NAND22 U62 ( .A(n363), .B(n360), .Q(n361) );
  NAND22 U63 ( .A(n363), .B(n360), .Q(n362) );
  NAND22 U64 ( .A(n363), .B(n360), .Q(n105) );
  INV3 U65 ( .A(Reset), .Q(n363) );
  INV3 U66 ( .A(n106), .Q(n360) );
  INV3 U67 ( .A(Din[5]), .Q(n390) );
  INV3 U68 ( .A(Din[3]), .Q(n393) );
  INV3 U69 ( .A(Din[1]), .Q(n394) );
  INV3 U70 ( .A(Din[2]), .Q(n392) );
  INV3 U71 ( .A(Din[0]), .Q(n395) );
  NOR20 U72 ( .A(Load), .B(Reset), .Q(n106) );
endmodule


module adder_40_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n50,
         n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n191, n194, n195, n196,
         n197, n198, n203, n204, n205, n206, n207, n208, n209, n212, n213,
         n214, n219, n220, n221, n222, n223, n224, n225, n226, n227, n230,
         n231, n232, n239, n240, n241, n242, n243, n244, n245, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n265, n266, n268, n269, n270, n271, n272, n273,
         n274, n275, n277, n278, n279, n280, n281, n547, n548, n549, n552,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U91 ( .A(n102), .B(n755), .C(n103), .Q(n101) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n755), .C(n141), .Q(n139) );
  OAI212 U159 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U165 ( .A(n158), .B(n755), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n760), .B(n755), .C(n756), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U189 ( .A(n176), .B(n755), .C(n177), .Q(n175) );
  OAI212 U201 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n778), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n776), .B(n778), .C(n774), .Q(n232) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n268), .B(n248), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  AOI212 U321 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  AOI212 U392 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U391 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  AOI212 U488 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U389 ( .A(n194), .B(n767), .C(n195), .Q(n191) );
  OAI212 U441 ( .A(n126), .B(n800), .C(n127), .Q(n123) );
  OAI212 U442 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  AOI212 U396 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U401 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U402 ( .A(n208), .B(n778), .C(n209), .Q(n207) );
  XNR22 U408 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U411 ( .A(n20), .B(n164), .Q(SUM[18]) );
  OAI212 U414 ( .A(n244), .B(n778), .C(n245), .Q(n243) );
  XNR22 U419 ( .A(n27), .B(n225), .Q(SUM[11]) );
  XNR22 U423 ( .A(n15), .B(n119), .Q(SUM[23]) );
  OAI212 U439 ( .A(n88), .B(n807), .C(n89), .Q(n85) );
  OAI212 U444 ( .A(n814), .B(n5), .C(n815), .Q(n56) );
  OAI212 U445 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U454 ( .A(n188), .B(n778), .C(n189), .Q(n187) );
  XNR22 U349 ( .A(n13), .B(n101), .Q(SUM[25]) );
  OAI212 U379 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  NOR24 U386 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR24 U387 ( .A(B[9]), .B(A[9]), .Q(n241) );
  OAI212 U388 ( .A(n129), .B(n755), .C(n130), .Q(n128) );
  OAI212 U416 ( .A(n755), .B(n91), .C(n92), .Q(n90) );
  XNR22 U427 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XNR22 U428 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XOR22 U433 ( .A(n22), .B(n755), .Q(SUM[16]) );
  XNR22 U435 ( .A(n21), .B(n175), .Q(SUM[17]) );
  XNR22 U436 ( .A(n24), .B(n196), .Q(SUM[14]) );
  XNR22 U443 ( .A(n26), .B(n214), .Q(SUM[12]) );
  AOI212 U363 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR24 U365 ( .A(B[15]), .B(A[15]), .Q(n185) );
  OAI212 U409 ( .A(n42), .B(n755), .C(n43), .Q(n41) );
  OAI212 U412 ( .A(n73), .B(n755), .C(n74), .Q(n72) );
  OAI212 U413 ( .A(n64), .B(n755), .C(n65), .Q(n63) );
  OAI212 U426 ( .A(n151), .B(n755), .C(n152), .Q(n146) );
  OAI212 U453 ( .A(n274), .B(n786), .C(n275), .Q(n273) );
  OAI212 U456 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U464 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  XNR22 U579 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NOR24 U617 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR22 U350 ( .A(n117), .B(n126), .Q(n115) );
  NAND20 U351 ( .A(n111), .B(n792), .Q(n73) );
  INV8 U352 ( .A(n247), .Q(n778) );
  AOI211 U353 ( .A(n769), .B(n203), .C(n204), .Q(n198) );
  NAND22 U354 ( .A(n761), .B(n122), .Q(n120) );
  INV2 U355 ( .A(n151), .Q(n761) );
  NOR20 U356 ( .A(n126), .B(n799), .Q(n122) );
  NOR22 U357 ( .A(n223), .B(n230), .Q(n221) );
  NOR23 U358 ( .A(B[11]), .B(A[11]), .Q(n223) );
  XNR22 U359 ( .A(n23), .B(n187), .Q(SUM[15]) );
  XNR22 U360 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U361 ( .A(n18), .B(n146), .Q(SUM[20]) );
  INV3 U362 ( .A(n204), .Q(n767) );
  INV6 U364 ( .A(n112), .Q(n752) );
  CLKIN6 U366 ( .A(n752), .Q(n753) );
  CLKIN8 U367 ( .A(n752), .Q(n754) );
  NAND23 U368 ( .A(n239), .B(n221), .Q(n219) );
  OAI211 U369 ( .A(n762), .B(n755), .C(n758), .Q(n108) );
  INV1 U370 ( .A(n111), .Q(n762) );
  XNR22 U371 ( .A(n243), .B(n29), .Q(SUM[9]) );
  NAND24 U372 ( .A(n171), .B(n153), .Q(n151) );
  NOR22 U373 ( .A(n185), .B(n194), .Q(n183) );
  AOI211 U374 ( .A(n754), .B(n820), .C(n819), .Q(n103) );
  NOR22 U375 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR22 U376 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NOR22 U377 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR22 U378 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR22 U380 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR23 U381 ( .A(B[13]), .B(A[13]), .Q(n205) );
  AOI211 U382 ( .A(n769), .B(n768), .C(n766), .Q(n209) );
  NOR21 U383 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NAND22 U384 ( .A(A[16]), .B(B[16]), .Q(n177) );
  XOR21 U385 ( .A(n33), .B(n262), .Q(SUM[5]) );
  XNR21 U390 ( .A(n28), .B(n232), .Q(SUM[10]) );
  OAI212 U393 ( .A(n120), .B(n755), .C(n121), .Q(n119) );
  CLKIN3 U394 ( .A(n145), .Q(n804) );
  NAND21 U395 ( .A(n805), .B(n145), .Q(n18) );
  AOI212 U397 ( .A(n754), .B(n84), .C(n85), .Q(n83) );
  NOR22 U398 ( .A(n181), .B(n219), .Q(n179) );
  CLKBU15 U399 ( .A(n178), .Q(n755) );
  INV1 U400 ( .A(n753), .Q(n758) );
  NAND21 U403 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NOR22 U404 ( .A(n260), .B(n265), .Q(n258) );
  INV2 U405 ( .A(n220), .Q(n769) );
  NOR24 U406 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR22 U407 ( .A(n271), .B(n274), .Q(n269) );
  OAI211 U410 ( .A(n197), .B(n778), .C(n198), .Q(n196) );
  NAND21 U415 ( .A(n111), .B(n790), .Q(n42) );
  AOI211 U417 ( .A(n754), .B(n97), .C(n98), .Q(n92) );
  NAND22 U418 ( .A(A[9]), .B(B[9]), .Q(n242) );
  INV1 U420 ( .A(n136), .Q(n800) );
  NAND21 U421 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND21 U422 ( .A(n111), .B(n820), .Q(n102) );
  NOR22 U424 ( .A(B[18]), .B(A[18]), .Q(n162) );
  XNR22 U425 ( .A(n11), .B(n81), .Q(SUM[27]) );
  OAI211 U429 ( .A(n82), .B(n755), .C(n83), .Q(n81) );
  AOI211 U430 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NAND20 U431 ( .A(n171), .B(n802), .Q(n158) );
  AOI211 U432 ( .A(n757), .B(n122), .C(n123), .Q(n121) );
  NOR21 U434 ( .A(n88), .B(n809), .Q(n84) );
  XNR22 U437 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR22 U438 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NOR24 U440 ( .A(n113), .B(n151), .Q(n111) );
  CLKIN2 U446 ( .A(n135), .Q(n799) );
  NAND22 U447 ( .A(A[10]), .B(B[10]), .Q(n231) );
  AOI210 U448 ( .A(n754), .B(n792), .C(n793), .Q(n74) );
  NAND21 U449 ( .A(n761), .B(n135), .Q(n129) );
  XOR20 U450 ( .A(n36), .B(n786), .Q(SUM[2]) );
  INV1 U451 ( .A(n277), .Q(n786) );
  XOR21 U452 ( .A(n778), .B(n30), .Q(SUM[8]) );
  AOI212 U455 ( .A(n784), .B(n781), .C(n782), .Q(n262) );
  INV2 U457 ( .A(n268), .Q(n784) );
  NAND21 U458 ( .A(n111), .B(n84), .Q(n82) );
  OAI211 U459 ( .A(n53), .B(n755), .C(n54), .Q(n52) );
  OAI210 U460 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  NOR22 U461 ( .A(n61), .B(n70), .Q(n59) );
  XNR22 U462 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U463 ( .A(n19), .B(n157), .Q(SUM[19]) );
  OAI212 U465 ( .A(n219), .B(n778), .C(n220), .Q(n214) );
  XNR21 U466 ( .A(n34), .B(n784), .Q(SUM[4]) );
  AOI212 U467 ( .A(n784), .B(n258), .C(n259), .Q(n257) );
  XOR22 U468 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NOR22 U469 ( .A(n241), .B(n244), .Q(n239) );
  NAND21 U470 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND21 U471 ( .A(n771), .B(n764), .Q(n188) );
  INV1 U472 ( .A(n5), .Q(n793) );
  NAND22 U473 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV2 U474 ( .A(n152), .Q(n757) );
  OAI210 U475 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  AOI210 U476 ( .A(n754), .B(n66), .C(n67), .Q(n65) );
  NAND21 U477 ( .A(n818), .B(n71), .Q(n10) );
  NAND21 U478 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NAND21 U479 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U480 ( .A(A[22]), .B(B[22]), .Q(n127) );
  INV3 U481 ( .A(n244), .Q(n775) );
  NAND20 U482 ( .A(n817), .B(n89), .Q(n12) );
  NAND20 U483 ( .A(n796), .B(n118), .Q(n15) );
  NAND20 U484 ( .A(n808), .B(n100), .Q(n13) );
  NAND20 U485 ( .A(n789), .B(n80), .Q(n11) );
  NAND20 U486 ( .A(n820), .B(n107), .Q(n14) );
  INV0 U487 ( .A(n106), .Q(n820) );
  INV0 U489 ( .A(n194), .Q(n765) );
  AOI210 U490 ( .A(n60), .B(n811), .C(n812), .Q(n47) );
  NOR21 U491 ( .A(n173), .B(n176), .Q(n171) );
  NAND22 U492 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U493 ( .A(B[1]), .B(A[1]), .Q(n279) );
  NOR23 U494 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND21 U495 ( .A(A[17]), .B(B[17]), .Q(n174) );
  INV1 U496 ( .A(n6), .Q(n792) );
  NOR20 U497 ( .A(n814), .B(n6), .Q(n55) );
  NAND20 U498 ( .A(n111), .B(n97), .Q(n91) );
  CLKIN0 U499 ( .A(n240), .Q(n774) );
  NOR22 U500 ( .A(n137), .B(n144), .Q(n135) );
  NOR22 U501 ( .A(n155), .B(n162), .Q(n153) );
  INV0 U502 ( .A(n137), .Q(n798) );
  NAND20 U503 ( .A(n779), .B(n256), .Q(n32) );
  INV1 U504 ( .A(n97), .Q(n809) );
  INV0 U505 ( .A(n88), .Q(n817) );
  NOR23 U506 ( .A(n205), .B(n212), .Q(n203) );
  INV0 U507 ( .A(n126), .Q(n797) );
  INV0 U508 ( .A(n99), .Q(n808) );
  INV0 U509 ( .A(n79), .Q(n789) );
  INV0 U510 ( .A(n70), .Q(n818) );
  INV0 U511 ( .A(n155), .Q(n801) );
  NAND20 U512 ( .A(n801), .B(n156), .Q(n19) );
  INV0 U513 ( .A(n163), .Q(n803) );
  NAND20 U514 ( .A(n59), .B(n811), .Q(n46) );
  NAND20 U515 ( .A(n768), .B(n213), .Q(n26) );
  XOR20 U516 ( .A(n281), .B(n37), .Q(SUM[1]) );
  CLKIN0 U517 ( .A(n278), .Q(n810) );
  NAND20 U518 ( .A(n775), .B(n245), .Q(n30) );
  NAND20 U519 ( .A(n783), .B(n275), .Q(n36) );
  INV0 U520 ( .A(n176), .Q(n759) );
  NAND20 U521 ( .A(n759), .B(n177), .Q(n22) );
  INV0 U522 ( .A(n117), .Q(n796) );
  INV0 U523 ( .A(n171), .Q(n760) );
  NAND20 U524 ( .A(n802), .B(n163), .Q(n20) );
  INV0 U525 ( .A(n213), .Q(n766) );
  INV0 U526 ( .A(n271), .Q(n806) );
  NAND20 U527 ( .A(n111), .B(n55), .Q(n53) );
  CLKIN0 U528 ( .A(n144), .Q(n805) );
  NOR20 U529 ( .A(n70), .B(n61), .Q(n549) );
  INV2 U530 ( .A(n548), .Q(n791) );
  NAND20 U531 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND21 U532 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NOR22 U533 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND21 U534 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND22 U535 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NOR22 U536 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR22 U537 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NAND20 U538 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U539 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND21 U540 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND21 U541 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND20 U542 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U543 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV3 U544 ( .A(n219), .Q(n771) );
  AOI210 U545 ( .A(n754), .B(n55), .C(n56), .Q(n54) );
  INV3 U546 ( .A(n60), .Q(n815) );
  NAND22 U547 ( .A(n97), .B(n77), .Q(n6) );
  AOI210 U548 ( .A(n757), .B(n135), .C(n136), .Q(n130) );
  INV3 U549 ( .A(n552), .Q(n764) );
  NAND22 U550 ( .A(n765), .B(n203), .Q(n552) );
  NAND20 U551 ( .A(n111), .B(n66), .Q(n64) );
  NAND22 U552 ( .A(n135), .B(n115), .Q(n113) );
  NAND22 U553 ( .A(n203), .B(n183), .Q(n181) );
  NAND22 U554 ( .A(n761), .B(n805), .Q(n140) );
  NAND22 U555 ( .A(n771), .B(n768), .Q(n208) );
  NAND22 U556 ( .A(n239), .B(n773), .Q(n226) );
  INV0 U557 ( .A(n172), .Q(n756) );
  INV3 U558 ( .A(n59), .Q(n814) );
  NAND22 U559 ( .A(n770), .B(n224), .Q(n27) );
  INV0 U560 ( .A(n223), .Q(n770) );
  NAND22 U561 ( .A(n797), .B(n127), .Q(n16) );
  NAND22 U562 ( .A(n258), .B(n250), .Q(n248) );
  NOR22 U563 ( .A(n252), .B(n255), .Q(n250) );
  NAND22 U564 ( .A(n794), .B(n174), .Q(n21) );
  INV3 U565 ( .A(n173), .Q(n794) );
  NAND22 U566 ( .A(n813), .B(n62), .Q(n9) );
  INV3 U567 ( .A(n61), .Q(n813) );
  NAND22 U568 ( .A(n798), .B(n138), .Q(n17) );
  NAND22 U569 ( .A(n795), .B(n242), .Q(n29) );
  INV0 U570 ( .A(n241), .Q(n795) );
  INV3 U571 ( .A(n107), .Q(n819) );
  INV0 U572 ( .A(n98), .Q(n807) );
  NAND22 U573 ( .A(n763), .B(n186), .Q(n23) );
  INV0 U574 ( .A(n185), .Q(n763) );
  NAND22 U575 ( .A(n788), .B(n206), .Q(n25) );
  INV0 U576 ( .A(n205), .Q(n788) );
  NOR21 U577 ( .A(n99), .B(n106), .Q(n97) );
  NAND22 U578 ( .A(n810), .B(n279), .Q(n37) );
  NAND22 U580 ( .A(n780), .B(n261), .Q(n33) );
  INV0 U581 ( .A(n260), .Q(n780) );
  INV0 U582 ( .A(n255), .Q(n779) );
  INV0 U583 ( .A(n274), .Q(n783) );
  INV3 U584 ( .A(n231), .Q(n772) );
  NAND22 U585 ( .A(n777), .B(n253), .Q(n31) );
  INV0 U586 ( .A(n252), .Q(n777) );
  XNR21 U587 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U588 ( .A(n806), .B(n272), .Q(n35) );
  NAND22 U589 ( .A(n765), .B(n195), .Q(n24) );
  NAND20 U590 ( .A(n771), .B(n203), .Q(n197) );
  XNR21 U591 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND22 U592 ( .A(n811), .B(n51), .Q(n8) );
  NAND22 U593 ( .A(n781), .B(n266), .Q(n34) );
  NAND22 U594 ( .A(n773), .B(n231), .Q(n28) );
  INV0 U595 ( .A(n239), .Q(n776) );
  AOI210 U596 ( .A(n754), .B(n790), .C(n45), .Q(n43) );
  NOR21 U597 ( .A(n70), .B(n6), .Q(n66) );
  NOR21 U598 ( .A(n79), .B(n88), .Q(n77) );
  AOI210 U599 ( .A(n172), .B(n802), .C(n803), .Q(n159) );
  AOI211 U600 ( .A(n757), .B(n805), .C(n804), .Q(n141) );
  AOI211 U601 ( .A(n769), .B(n764), .C(n191), .Q(n189) );
  NAND20 U602 ( .A(n792), .B(n811), .Q(n548) );
  INV3 U603 ( .A(n162), .Q(n802) );
  INV3 U604 ( .A(n212), .Q(n768) );
  INV3 U605 ( .A(n230), .Q(n773) );
  INV3 U606 ( .A(n265), .Q(n781) );
  INV3 U607 ( .A(n547), .Q(n790) );
  NAND22 U608 ( .A(n549), .B(n791), .Q(n547) );
  INV3 U609 ( .A(n266), .Q(n782) );
  INV3 U610 ( .A(n51), .Q(n812) );
  NOR21 U611 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR22 U612 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR21 U613 ( .A(B[29]), .B(A[29]), .Q(n61) );
  XNR21 U614 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U615 ( .A(n816), .B(n40), .Q(n7) );
  NAND22 U616 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR22 U618 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR22 U619 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR22 U620 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR22 U621 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR22 U622 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR22 U623 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR21 U624 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR23 U625 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND22 U626 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND21 U627 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND22 U628 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND22 U629 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND22 U630 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U631 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND21 U632 ( .A(A[13]), .B(B[13]), .Q(n206) );
  INV3 U633 ( .A(n38), .Q(SUM[0]) );
  NAND20 U634 ( .A(n787), .B(n281), .Q(n38) );
  INV3 U635 ( .A(n280), .Q(n787) );
  NOR20 U636 ( .A(B[0]), .B(A[0]), .Q(n280) );
  INV3 U637 ( .A(n50), .Q(n811) );
  NOR21 U638 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND22 U639 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U640 ( .A(n39), .Q(n816) );
  NOR21 U641 ( .A(B[31]), .B(A[31]), .Q(n39) );
  AOI210 U642 ( .A(n240), .B(n773), .C(n772), .Q(n227) );
endmodule


module adder_40 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_40_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_39_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n427, n579, n726,
         n729, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n871;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  AOI212 U195 ( .A(n179), .B(n247), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U483 ( .A(n99), .B(n107), .C(n100), .Q(n98) );
  OAI212 U510 ( .A(n79), .B(n89), .C(n80), .Q(n78) );
  AOI212 U529 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  OAI212 U475 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  AOI212 U458 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI212 U481 ( .A(n803), .B(n91), .C(n92), .Q(n90) );
  OAI212 U467 ( .A(n274), .B(n869), .C(n275), .Q(n273) );
  OAI212 U511 ( .A(n129), .B(n803), .C(n130), .Q(n128) );
  OAI212 U514 ( .A(n158), .B(n803), .C(n159), .Q(n157) );
  OAI212 U369 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U512 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U652 ( .A(n819), .B(n806), .C(n816), .Q(n579) );
  XNR22 U406 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U407 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U420 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NOR24 U441 ( .A(B[26]), .B(A[26]), .Q(n88) );
  OAI212 U442 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U464 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  AOI212 U465 ( .A(n805), .B(n822), .C(n825), .Q(n103) );
  NOR24 U468 ( .A(B[22]), .B(A[22]), .Q(n126) );
  OAI212 U505 ( .A(n82), .B(n803), .C(n83), .Q(n81) );
  OAI212 U513 ( .A(n155), .B(n163), .C(n156), .Q(n154) );
  NOR24 U360 ( .A(B[21]), .B(A[21]), .Q(n137) );
  OAI212 U382 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U414 ( .A(n860), .B(n188), .C(n189), .Q(n187) );
  NAND28 U356 ( .A(n812), .B(n842), .Q(n726) );
  OAI212 U412 ( .A(n194), .B(n847), .C(n195), .Q(n191) );
  OAI212 U418 ( .A(n860), .B(n219), .C(n220), .Q(n214) );
  OAI212 U435 ( .A(n226), .B(n860), .C(n227), .Q(n225) );
  OAI212 U436 ( .A(n208), .B(n860), .C(n209), .Q(n207) );
  OAI212 U437 ( .A(n857), .B(n860), .C(n855), .Q(n232) );
  OAI212 U438 ( .A(n197), .B(n860), .C(n198), .Q(n196) );
  OAI212 U444 ( .A(n140), .B(n802), .C(n141), .Q(n139) );
  OAI212 U445 ( .A(n808), .B(n802), .C(n804), .Q(n164) );
  INV2 U349 ( .A(n172), .Q(n804) );
  INV3 U350 ( .A(n135), .Q(n818) );
  OAI212 U351 ( .A(n176), .B(n802), .C(n177), .Q(n175) );
  CLKIN15 U352 ( .A(n801), .Q(n802) );
  NOR23 U353 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR24 U354 ( .A(B[19]), .B(A[19]), .Q(n155) );
  INV6 U355 ( .A(n152), .Q(n806) );
  NAND24 U357 ( .A(n427), .B(n43), .Q(n41) );
  INV1 U358 ( .A(n274), .Q(n866) );
  OAI210 U359 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  AOI211 U361 ( .A(n865), .B(n258), .C(n259), .Q(n257) );
  NOR24 U362 ( .A(n155), .B(n162), .Q(n153) );
  OAI212 U363 ( .A(n810), .B(n803), .C(n729), .Q(n108) );
  INV10 U364 ( .A(n801), .Q(n803) );
  INV1 U365 ( .A(n111), .Q(n810) );
  NOR24 U366 ( .A(B[25]), .B(A[25]), .Q(n99) );
  OAI212 U367 ( .A(n151), .B(n802), .C(n152), .Q(n146) );
  NOR24 U368 ( .A(n79), .B(n88), .Q(n77) );
  NOR22 U370 ( .A(B[24]), .B(A[24]), .Q(n106) );
  OAI211 U371 ( .A(n88), .B(n826), .C(n89), .Q(n85) );
  INV1 U372 ( .A(n98), .Q(n826) );
  OAI211 U373 ( .A(n5), .B(n70), .C(n71), .Q(n67) );
  NAND22 U374 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND22 U375 ( .A(A[26]), .B(B[26]), .Q(n89) );
  INV1 U376 ( .A(n106), .Q(n822) );
  NOR23 U377 ( .A(n830), .B(n6), .Q(n55) );
  NOR22 U378 ( .A(A[12]), .B(B[12]), .Q(n212) );
  NAND24 U379 ( .A(n171), .B(n153), .Q(n151) );
  NAND23 U380 ( .A(n239), .B(n221), .Q(n219) );
  NOR22 U381 ( .A(n223), .B(n230), .Q(n221) );
  OAI211 U383 ( .A(n244), .B(n860), .C(n245), .Q(n243) );
  INV0 U384 ( .A(n244), .Q(n856) );
  NOR22 U385 ( .A(n241), .B(n244), .Q(n239) );
  NOR22 U386 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR22 U387 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR22 U388 ( .A(n260), .B(n265), .Q(n258) );
  NOR22 U389 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR22 U390 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR22 U391 ( .A(B[16]), .B(A[16]), .Q(n176) );
  INV6 U392 ( .A(n178), .Q(n801) );
  NOR23 U393 ( .A(n181), .B(n219), .Q(n179) );
  NAND24 U394 ( .A(A[16]), .B(B[16]), .Q(n177) );
  AOI211 U395 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND23 U396 ( .A(n203), .B(n183), .Q(n181) );
  NOR23 U397 ( .A(B[27]), .B(A[27]), .Q(n79) );
  INV3 U398 ( .A(n114), .Q(n816) );
  INV3 U399 ( .A(n113), .Q(n819) );
  NOR23 U400 ( .A(n137), .B(n144), .Q(n135) );
  NOR23 U401 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR22 U402 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR22 U403 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR22 U404 ( .A(n173), .B(n176), .Q(n171) );
  NOR22 U405 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NOR21 U408 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND22 U409 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U410 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR23 U411 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR22 U413 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NOR22 U415 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR23 U416 ( .A(n205), .B(n212), .Q(n203) );
  NOR23 U417 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND22 U419 ( .A(n111), .B(n824), .Q(n73) );
  NOR21 U421 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U422 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND22 U423 ( .A(A[8]), .B(B[8]), .Q(n245) );
  XNR21 U424 ( .A(n21), .B(n175), .Q(SUM[17]) );
  INV2 U425 ( .A(n804), .Q(n800) );
  NAND24 U426 ( .A(n726), .B(n103), .Q(n101) );
  NAND22 U427 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND22 U428 ( .A(n809), .B(n122), .Q(n120) );
  NAND21 U429 ( .A(n111), .B(n822), .Q(n102) );
  AOI211 U430 ( .A(n806), .B(n122), .C(n123), .Q(n121) );
  OAI211 U431 ( .A(n126), .B(n815), .C(n127), .Q(n123) );
  AOI212 U432 ( .A(n805), .B(n97), .C(n98), .Q(n92) );
  OAI212 U433 ( .A(n120), .B(n803), .C(n121), .Q(n119) );
  INV3 U434 ( .A(n247), .Q(n860) );
  OAI211 U439 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  INV1 U440 ( .A(n220), .Q(n852) );
  NAND24 U443 ( .A(n135), .B(n115), .Q(n113) );
  AOI212 U446 ( .A(n805), .B(n55), .C(n56), .Q(n54) );
  INV1 U447 ( .A(n136), .Q(n815) );
  NOR23 U448 ( .A(n61), .B(n70), .Q(n59) );
  INV2 U449 ( .A(n70), .Q(n833) );
  NOR22 U450 ( .A(n70), .B(n6), .Q(n66) );
  NAND22 U451 ( .A(n111), .B(n55), .Q(n53) );
  NOR23 U452 ( .A(B[28]), .B(A[28]), .Q(n70) );
  AOI212 U453 ( .A(n805), .B(n84), .C(n85), .Q(n83) );
  XNR22 U454 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NAND22 U455 ( .A(B[17]), .B(A[17]), .Q(n174) );
  AOI212 U456 ( .A(n805), .B(n44), .C(n45), .Q(n43) );
  XNR22 U457 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NAND22 U459 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NOR21 U460 ( .A(n126), .B(n818), .Q(n122) );
  CLKIN3 U461 ( .A(n107), .Q(n825) );
  OAI211 U462 ( .A(n5), .B(n830), .C(n828), .Q(n56) );
  OAI211 U463 ( .A(n5), .B(n46), .C(n47), .Q(n45) );
  INV1 U466 ( .A(n5), .Q(n827) );
  OAI212 U469 ( .A(n64), .B(n803), .C(n65), .Q(n63) );
  XNR22 U470 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND21 U471 ( .A(A[30]), .B(B[30]), .Q(n51) );
  OAI212 U472 ( .A(n73), .B(n803), .C(n74), .Q(n72) );
  AOI212 U473 ( .A(n805), .B(n824), .C(n827), .Q(n74) );
  NAND21 U474 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND22 U476 ( .A(B[19]), .B(A[19]), .Q(n156) );
  XNR22 U477 ( .A(n8), .B(n52), .Q(SUM[30]) );
  OAI212 U478 ( .A(n53), .B(n803), .C(n54), .Q(n52) );
  NOR22 U479 ( .A(n46), .B(n6), .Q(n44) );
  INV2 U480 ( .A(n97), .Q(n823) );
  NOR23 U482 ( .A(n99), .B(n106), .Q(n97) );
  INV6 U484 ( .A(n579), .Q(n805) );
  OAI212 U485 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NAND22 U486 ( .A(B[22]), .B(A[22]), .Q(n127) );
  NOR21 U487 ( .A(n88), .B(n823), .Q(n84) );
  NAND24 U488 ( .A(n97), .B(n77), .Q(n6) );
  AOI212 U489 ( .A(n805), .B(n66), .C(n67), .Q(n65) );
  NOR23 U490 ( .A(n185), .B(n194), .Q(n183) );
  NAND22 U491 ( .A(n111), .B(n44), .Q(n42) );
  NAND21 U492 ( .A(n111), .B(n66), .Q(n64) );
  NAND22 U493 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NOR24 U494 ( .A(n113), .B(n151), .Q(n111) );
  NAND21 U495 ( .A(n851), .B(n190), .Q(n188) );
  AOI210 U496 ( .A(n852), .B(n190), .C(n191), .Q(n189) );
  NOR24 U497 ( .A(B[17]), .B(A[17]), .Q(n173) );
  INV2 U498 ( .A(n59), .Q(n830) );
  NAND24 U499 ( .A(n811), .B(n842), .Q(n427) );
  NAND21 U500 ( .A(n111), .B(n84), .Q(n82) );
  NAND21 U501 ( .A(A[23]), .B(B[23]), .Q(n118) );
  INV6 U502 ( .A(n802), .Q(n842) );
  AOI211 U503 ( .A(n60), .B(n837), .C(n836), .Q(n47) );
  INV0 U504 ( .A(n162), .Q(n814) );
  NOR22 U506 ( .A(n271), .B(n274), .Q(n269) );
  INV0 U507 ( .A(n213), .Q(n849) );
  NAND22 U508 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND22 U509 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NOR21 U515 ( .A(B[1]), .B(A[1]), .Q(n278) );
  INV2 U516 ( .A(n102), .Q(n812) );
  NAND20 U517 ( .A(n111), .B(n97), .Q(n91) );
  CLKIN0 U518 ( .A(n171), .Q(n808) );
  NOR24 U519 ( .A(n117), .B(n126), .Q(n115) );
  NOR24 U520 ( .A(n252), .B(n255), .Q(n250) );
  AOI212 U521 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  INV0 U522 ( .A(n144), .Q(n838) );
  INV0 U523 ( .A(n230), .Q(n853) );
  AOI210 U524 ( .A(n865), .B(n863), .C(n864), .Q(n262) );
  INV0 U525 ( .A(n266), .Q(n864) );
  NOR20 U526 ( .A(n194), .B(n846), .Q(n190) );
  NAND21 U527 ( .A(n851), .B(n848), .Q(n208) );
  CLKIN0 U528 ( .A(n204), .Q(n847) );
  INV0 U530 ( .A(n212), .Q(n848) );
  INV0 U531 ( .A(n265), .Q(n863) );
  INV0 U532 ( .A(n277), .Q(n869) );
  INV0 U533 ( .A(n271), .Q(n867) );
  NOR22 U534 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND22 U535 ( .A(B[14]), .B(A[14]), .Q(n195) );
  NAND22 U536 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND24 U537 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND21 U538 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U539 ( .A(B[3]), .B(A[3]), .Q(n272) );
  NAND20 U540 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND22 U541 ( .A(A[12]), .B(B[12]), .Q(n213) );
  XOR21 U542 ( .A(n30), .B(n860), .Q(SUM[8]) );
  XNR20 U543 ( .A(n34), .B(n865), .Q(SUM[4]) );
  NAND20 U544 ( .A(n866), .B(n275), .Q(n36) );
  NAND20 U545 ( .A(n868), .B(n279), .Q(n37) );
  XOR20 U546 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND20 U547 ( .A(n867), .B(n272), .Q(n35) );
  NAND20 U548 ( .A(n871), .B(n281), .Q(n38) );
  INV3 U549 ( .A(n6), .Q(n824) );
  INV3 U550 ( .A(n42), .Q(n811) );
  INV3 U551 ( .A(n151), .Q(n809) );
  INV3 U552 ( .A(n219), .Q(n851) );
  AOI210 U553 ( .A(n819), .B(n806), .C(n816), .Q(n729) );
  NAND20 U554 ( .A(n809), .B(n135), .Q(n129) );
  INV3 U555 ( .A(n60), .Q(n828) );
  NAND22 U556 ( .A(n851), .B(n203), .Q(n197) );
  AOI210 U557 ( .A(n852), .B(n203), .C(n204), .Q(n198) );
  INV3 U558 ( .A(n239), .Q(n857) );
  INV0 U559 ( .A(n240), .Q(n855) );
  INV3 U560 ( .A(n268), .Q(n865) );
  INV3 U561 ( .A(n203), .Q(n846) );
  NAND20 U562 ( .A(n171), .B(n814), .Q(n158) );
  AOI210 U563 ( .A(n800), .B(n814), .C(n813), .Q(n159) );
  INV3 U564 ( .A(n163), .Q(n813) );
  NAND20 U565 ( .A(n809), .B(n838), .Q(n140) );
  AOI210 U566 ( .A(n806), .B(n838), .C(n839), .Q(n141) );
  INV3 U567 ( .A(n145), .Q(n839) );
  AOI210 U568 ( .A(n852), .B(n848), .C(n849), .Q(n209) );
  NAND20 U569 ( .A(n239), .B(n853), .Q(n226) );
  AOI210 U570 ( .A(n240), .B(n853), .C(n854), .Q(n227) );
  INV3 U571 ( .A(n231), .Q(n854) );
  INV3 U572 ( .A(n51), .Q(n836) );
  NAND22 U573 ( .A(n59), .B(n837), .Q(n46) );
  INV0 U574 ( .A(n155), .Q(n840) );
  INV0 U575 ( .A(n126), .Q(n821) );
  INV0 U576 ( .A(n194), .Q(n844) );
  INV0 U577 ( .A(n88), .Q(n831) );
  INV0 U578 ( .A(n137), .Q(n817) );
  INV0 U579 ( .A(n260), .Q(n862) );
  INV0 U580 ( .A(n255), .Q(n861) );
  INV0 U581 ( .A(n176), .Q(n807) );
  INV0 U582 ( .A(n99), .Q(n832) );
  INV0 U583 ( .A(n79), .Q(n835) );
  INV0 U584 ( .A(n117), .Q(n820) );
  INV0 U585 ( .A(n205), .Q(n845) );
  INV0 U586 ( .A(n185), .Q(n843) );
  INV3 U587 ( .A(n61), .Q(n829) );
  INV0 U588 ( .A(n241), .Q(n858) );
  INV0 U589 ( .A(n252), .Q(n859) );
  INV0 U590 ( .A(n223), .Q(n850) );
  INV3 U591 ( .A(n173), .Q(n841) );
  INV3 U592 ( .A(n278), .Q(n868) );
  NOR21 U593 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U594 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NAND22 U595 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U596 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND21 U597 ( .A(B[9]), .B(A[9]), .Q(n242) );
  NAND21 U598 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND21 U599 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND21 U600 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND21 U601 ( .A(B[11]), .B(A[11]), .Q(n224) );
  INV3 U602 ( .A(n50), .Q(n837) );
  NOR21 U603 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND22 U604 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND22 U605 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV3 U606 ( .A(n39), .Q(n834) );
  INV3 U607 ( .A(n280), .Q(n871) );
  NOR21 U608 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U609 ( .A(n832), .B(n100), .Q(n13) );
  NAND20 U610 ( .A(n831), .B(n89), .Q(n12) );
  NAND20 U611 ( .A(n829), .B(n62), .Q(n9) );
  NAND20 U612 ( .A(n833), .B(n71), .Q(n10) );
  XNR21 U613 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U614 ( .A(n156), .B(n840), .Q(n19) );
  XNR21 U615 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND20 U616 ( .A(n821), .B(n127), .Q(n16) );
  XNR21 U617 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND20 U618 ( .A(n820), .B(n118), .Q(n15) );
  NAND20 U619 ( .A(n841), .B(n174), .Q(n21) );
  XNR21 U620 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND20 U621 ( .A(n838), .B(n145), .Q(n18) );
  NAND22 U622 ( .A(n834), .B(n40), .Q(n7) );
  NAND20 U623 ( .A(n835), .B(n80), .Q(n11) );
  NAND20 U624 ( .A(n837), .B(n51), .Q(n8) );
  XNR21 U625 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND20 U626 ( .A(n822), .B(n107), .Q(n14) );
  XNR21 U627 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND20 U628 ( .A(n163), .B(n814), .Q(n20) );
  XNR21 U629 ( .A(n17), .B(n139), .Q(SUM[21]) );
  NAND20 U630 ( .A(n817), .B(n138), .Q(n17) );
  XNR21 U631 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U632 ( .A(n859), .B(n253), .Q(n31) );
  XOR20 U633 ( .A(n22), .B(n802), .Q(SUM[16]) );
  NAND20 U634 ( .A(n807), .B(n177), .Q(n22) );
  XNR21 U635 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U636 ( .A(n844), .B(n195), .Q(n24) );
  XNR21 U637 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U638 ( .A(n845), .B(n206), .Q(n25) );
  XNR21 U639 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U640 ( .A(n853), .B(n231), .Q(n28) );
  XNR21 U641 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U642 ( .A(n850), .B(n224), .Q(n27) );
  NAND20 U643 ( .A(n856), .B(n245), .Q(n30) );
  NAND20 U644 ( .A(n863), .B(n266), .Q(n34) );
  XOR21 U645 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND20 U646 ( .A(n862), .B(n261), .Q(n33) );
  XNR21 U647 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U648 ( .A(n843), .B(n186), .Q(n23) );
  XNR21 U649 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U650 ( .A(n858), .B(n242), .Q(n29) );
  XNR21 U651 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U653 ( .A(n848), .B(n213), .Q(n26) );
  XOR21 U654 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND20 U655 ( .A(n861), .B(n256), .Q(n32) );
  XNR21 U656 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XOR21 U657 ( .A(n36), .B(n869), .Q(SUM[2]) );
  INV3 U658 ( .A(n38), .Q(SUM[0]) );
  AOI210 U659 ( .A(n806), .B(n135), .C(n136), .Q(n130) );
endmodule


module adder_39 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_39_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module reg_11 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31,
         n34, n50, n52, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n54, n55, n56, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n108, n109, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393;

  DF3 Dout_reg_19_ ( .D(n69), .C(Clk), .Q(Dout[19]), .QN(n13) );
  DF3 Dout_reg_18_ ( .D(n70), .C(Clk), .Q(Dout[18]), .QN(n11) );
  DF3 Dout_reg_16_ ( .D(n72), .C(Clk), .Q(Dout[16]), .QN(n7) );
  DF3 Dout_reg_15_ ( .D(n73), .C(Clk), .Q(Dout[15]), .QN(n5) );
  DF3 Dout_reg_14_ ( .D(n86), .C(Clk), .Q(Dout[14]), .QN(n56) );
  DF3 Dout_reg_12_ ( .D(n88), .C(Clk), .Q(Dout[12]), .QN(n79) );
  DF3 Dout_reg_11_ ( .D(n89), .C(Clk), .Q(Dout[11]), .QN(n55) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n78) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n77) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n76) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n75) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n74) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n84) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n83) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n81) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n80) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n85) );
  DF3 Dout_reg_17_ ( .D(n71), .C(Clk), .Q(Dout[17]), .QN(n9) );
  DF3 Dout_reg_23_ ( .D(n65), .C(Clk), .Q(Dout[23]), .QN(n21) );
  DF3 Dout_reg_13_ ( .D(n87), .C(Clk), .Q(Dout[13]), .QN(n54) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n82) );
  DF3 Dout_reg_29_ ( .D(n59), .C(Clk), .Q(Dout[29]), .QN(n34) );
  DF3 Dout_reg_27_ ( .D(n61), .C(Clk), .Q(Dout[27]), .QN(n29) );
  OAI222 U3 ( .A(n80), .B(n358), .C(n360), .D(n391), .Q(n99) );
  OAI222 U4 ( .A(n81), .B(n358), .C(n359), .D(n392), .Q(n98) );
  OAI222 U5 ( .A(n82), .B(n358), .C(n108), .D(n393), .Q(n97) );
  OAI222 U6 ( .A(n83), .B(n358), .C(n360), .D(n389), .Q(n96) );
  OAI222 U7 ( .A(n84), .B(n358), .C(n359), .D(n381), .Q(n95) );
  OAI222 U8 ( .A(n74), .B(n358), .C(n108), .D(n380), .Q(n94) );
  OAI222 U9 ( .A(n75), .B(n358), .C(n360), .D(n383), .Q(n93) );
  OAI222 U10 ( .A(n76), .B(n358), .C(n359), .D(n382), .Q(n92) );
  OAI222 U11 ( .A(n77), .B(n358), .C(n108), .D(n387), .Q(n91) );
  OAI222 U12 ( .A(n78), .B(n358), .C(n360), .D(n388), .Q(n90) );
  OAI222 U13 ( .A(n55), .B(n358), .C(n359), .D(n385), .Q(n89) );
  OAI222 U14 ( .A(n79), .B(n358), .C(n108), .D(n386), .Q(n88) );
  OAI222 U15 ( .A(n54), .B(n358), .C(n360), .D(n384), .Q(n87) );
  OAI222 U16 ( .A(n56), .B(n358), .C(n359), .D(n379), .Q(n86) );
  OAI222 U17 ( .A(n5), .B(n358), .C(n108), .D(n378), .Q(n73) );
  OAI222 U18 ( .A(n7), .B(n358), .C(n360), .D(n377), .Q(n72) );
  OAI222 U19 ( .A(n9), .B(n358), .C(n359), .D(n375), .Q(n71) );
  OAI222 U20 ( .A(n11), .B(n358), .C(n108), .D(n374), .Q(n70) );
  OAI222 U21 ( .A(n13), .B(n358), .C(n360), .D(n376), .Q(n69) );
  OAI222 U22 ( .A(n15), .B(n358), .C(n359), .D(n373), .Q(n68) );
  OAI222 U23 ( .A(n17), .B(n358), .C(n108), .D(n372), .Q(n67) );
  OAI222 U24 ( .A(n19), .B(n358), .C(n360), .D(n371), .Q(n66) );
  OAI222 U25 ( .A(n21), .B(n358), .C(n359), .D(n370), .Q(n65) );
  OAI222 U26 ( .A(n23), .B(n358), .C(n108), .D(n369), .Q(n64) );
  OAI222 U27 ( .A(n25), .B(n358), .C(n360), .D(n368), .Q(n63) );
  OAI222 U28 ( .A(n27), .B(n358), .C(n359), .D(n367), .Q(n62) );
  OAI222 U29 ( .A(n29), .B(n358), .C(n366), .D(n108), .Q(n61) );
  OAI222 U30 ( .A(n31), .B(n358), .C(n360), .D(n365), .Q(n60) );
  OAI222 U31 ( .A(n34), .B(n358), .C(n359), .D(n364), .Q(n59) );
  OAI222 U32 ( .A(n50), .B(n358), .C(n363), .D(n108), .Q(n58) );
  OAI222 U33 ( .A(n52), .B(n358), .C(n362), .D(n360), .Q(n57) );
  OAI222 U34 ( .A(n85), .B(n358), .C(n359), .D(n390), .Q(n100) );
  DF1 Dout_reg_31_ ( .D(n57), .C(Clk), .Q(Dout[31]), .QN(n52) );
  DF1 Dout_reg_28_ ( .D(n60), .C(Clk), .Q(Dout[28]), .QN(n31) );
  DF1 Dout_reg_26_ ( .D(n62), .C(Clk), .Q(Dout[26]), .QN(n27) );
  DF1 Dout_reg_20_ ( .D(n68), .C(Clk), .Q(Dout[20]), .QN(n15) );
  DF1 Dout_reg_25_ ( .D(n63), .C(Clk), .Q(Dout[25]), .QN(n25) );
  DF1 Dout_reg_24_ ( .D(n64), .C(Clk), .Q(Dout[24]), .QN(n23) );
  DF1 Dout_reg_22_ ( .D(n66), .C(Clk), .Q(Dout[22]), .QN(n19) );
  DF1 Dout_reg_30_ ( .D(n58), .C(Clk), .Q(Dout[30]), .QN(n50) );
  DF3 Dout_reg_21_ ( .D(n67), .C(Clk), .Q(Dout[21]), .QN(n17) );
  INV3 U35 ( .A(Din[31]), .Q(n362) );
  INV3 U36 ( .A(Din[28]), .Q(n365) );
  INV3 U37 ( .A(Din[30]), .Q(n363) );
  INV3 U38 ( .A(Din[29]), .Q(n364) );
  INV2 U39 ( .A(Din[27]), .Q(n366) );
  INV3 U40 ( .A(Din[18]), .Q(n374) );
  INV2 U41 ( .A(Din[16]), .Q(n377) );
  CLKIN3 U42 ( .A(Din[15]), .Q(n378) );
  INV2 U43 ( .A(Din[14]), .Q(n379) );
  INV2 U44 ( .A(Din[26]), .Q(n367) );
  INV2 U45 ( .A(Din[25]), .Q(n368) );
  INV2 U46 ( .A(Din[22]), .Q(n371) );
  INV2 U47 ( .A(Din[20]), .Q(n373) );
  INV2 U48 ( .A(Din[23]), .Q(n370) );
  INV2 U49 ( .A(Din[19]), .Q(n376) );
  INV2 U50 ( .A(Din[17]), .Q(n375) );
  INV2 U51 ( .A(Din[24]), .Q(n369) );
  INV2 U52 ( .A(Din[21]), .Q(n372) );
  CLKIN3 U53 ( .A(Din[9]), .Q(n387) );
  NAND22 U54 ( .A(n361), .B(n358), .Q(n359) );
  NAND22 U55 ( .A(n361), .B(n358), .Q(n360) );
  NAND22 U56 ( .A(n361), .B(n358), .Q(n108) );
  INV3 U57 ( .A(Reset), .Q(n361) );
  INV3 U58 ( .A(n109), .Q(n358) );
  INV3 U59 ( .A(Din[13]), .Q(n384) );
  INV3 U60 ( .A(Din[10]), .Q(n388) );
  INV3 U61 ( .A(Din[11]), .Q(n385) );
  INV3 U62 ( .A(Din[7]), .Q(n383) );
  INV3 U63 ( .A(Din[8]), .Q(n382) );
  INV3 U64 ( .A(Din[12]), .Q(n386) );
  INV3 U65 ( .A(Din[3]), .Q(n393) );
  INV3 U66 ( .A(Din[6]), .Q(n380) );
  INV3 U67 ( .A(Din[1]), .Q(n391) );
  INV3 U68 ( .A(Din[2]), .Q(n392) );
  INV3 U69 ( .A(Din[4]), .Q(n389) );
  INV3 U70 ( .A(Din[5]), .Q(n381) );
  INV3 U71 ( .A(Din[0]), .Q(n390) );
  NOR20 U72 ( .A(Load), .B(Reset), .Q(n109) );
endmodule


module reg_10 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n4, n6, n8, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n53, n54, n55, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n104, n17, n19, n21, n23, n25, n27,
         n29, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n101, n102, n103, n105, n106,
         n107, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325;

  DF3 Dout_reg_16_ ( .D(n71), .C(Clk), .Q(Dout[16]), .QN(n4) );
  DF3 Dout_reg_15_ ( .D(n85), .C(Clk), .Q(Dout[15]), .QN(n72) );
  DF3 Dout_reg_14_ ( .D(n86), .C(Clk), .Q(Dout[14]), .QN(n55) );
  DF3 Dout_reg_13_ ( .D(n87), .C(Clk), .Q(Dout[13]), .QN(n54) );
  DF3 Dout_reg_12_ ( .D(n88), .C(Clk), .Q(Dout[12]), .QN(n53) );
  DF3 Dout_reg_11_ ( .D(n89), .C(Clk), .Q(Dout[11]), .QN(n77) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n76) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n74) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n73) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n78) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n82) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n81) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n84) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n83) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n75) );
  DF3 Dout_reg_19_ ( .D(n68), .C(Clk), .Q(Dout[19]) );
  DF3 Dout_reg_18_ ( .D(n69), .C(Clk), .Q(Dout[18]), .QN(n8) );
  DF3 Dout_reg_17_ ( .D(n70), .C(Clk), .Q(Dout[17]), .QN(n6) );
  DF3 Dout_reg_23_ ( .D(n64), .C(Clk), .Q(Dout[23]), .QN(n18) );
  DF3 Dout_reg_21_ ( .D(n66), .C(Clk), .Q(Dout[21]), .QN(n14) );
  DF3 Dout_reg_22_ ( .D(n65), .C(Clk), .Q(Dout[22]), .QN(n16) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n79) );
  DF3 Dout_reg_20_ ( .D(n67), .C(Clk), .Q(Dout[20]), .QN(n12) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n80) );
  DF3 Dout_reg_24_ ( .D(n63), .C(Clk), .Q(Dout[24]), .QN(n20) );
  OAI212 U3 ( .A(n84), .B(n321), .C(n17), .Q(n99) );
  OAI212 U5 ( .A(n79), .B(n321), .C(n21), .Q(n98) );
  OAI212 U7 ( .A(n80), .B(n321), .C(n23), .Q(n97) );
  OAI212 U9 ( .A(n81), .B(n321), .C(n25), .Q(n96) );
  OAI212 U11 ( .A(n82), .B(n321), .C(n27), .Q(n95) );
  OAI212 U13 ( .A(n78), .B(n321), .C(n29), .Q(n94) );
  OAI212 U15 ( .A(n73), .B(n321), .C(n31), .Q(n93) );
  OAI212 U17 ( .A(n74), .B(n321), .C(n33), .Q(n92) );
  OAI212 U19 ( .A(n75), .B(n321), .C(n34), .Q(n91) );
  OAI212 U21 ( .A(n76), .B(n321), .C(n35), .Q(n90) );
  OAI212 U23 ( .A(n77), .B(n321), .C(n36), .Q(n89) );
  OAI212 U25 ( .A(n53), .B(n321), .C(n37), .Q(n88) );
  OAI212 U27 ( .A(n54), .B(n321), .C(n38), .Q(n87) );
  OAI212 U29 ( .A(n55), .B(n321), .C(n39), .Q(n86) );
  OAI212 U31 ( .A(n72), .B(n321), .C(n40), .Q(n85) );
  OAI212 U33 ( .A(n4), .B(n321), .C(n41), .Q(n71) );
  OAI212 U35 ( .A(n6), .B(n321), .C(n42), .Q(n70) );
  OAI212 U37 ( .A(n8), .B(n321), .C(n43), .Q(n69) );
  OAI212 U41 ( .A(n12), .B(n321), .C(n45), .Q(n67) );
  OAI212 U43 ( .A(n14), .B(n321), .C(n46), .Q(n66) );
  OAI212 U45 ( .A(n16), .B(n321), .C(n47), .Q(n65) );
  OAI212 U47 ( .A(n18), .B(n321), .C(n48), .Q(n64) );
  OAI212 U49 ( .A(n20), .B(n321), .C(n49), .Q(n63) );
  OAI212 U51 ( .A(n22), .B(n321), .C(n50), .Q(n62) );
  OAI212 U53 ( .A(n24), .B(n321), .C(n51), .Q(n61) );
  OAI212 U55 ( .A(n26), .B(n321), .C(n52), .Q(n60) );
  OAI212 U57 ( .A(n28), .B(n321), .C(n101), .Q(n59) );
  OAI212 U59 ( .A(n30), .B(n321), .C(n102), .Q(n58) );
  OAI212 U61 ( .A(n32), .B(n321), .C(n103), .Q(n57) );
  OAI212 U63 ( .A(n104), .B(n321), .C(n105), .Q(n56) );
  OAI212 U65 ( .A(n83), .B(n321), .C(n106), .Q(n100) );
  DF1 Dout_reg_30_ ( .D(n57), .C(Clk), .Q(Dout[30]), .QN(n32) );
  DF1 Dout_reg_29_ ( .D(n58), .C(Clk), .Q(Dout[29]), .QN(n30) );
  DF1 Dout_reg_28_ ( .D(n59), .C(Clk), .Q(Dout[28]), .QN(n28) );
  DF1 Dout_reg_31_ ( .D(n56), .C(Clk), .Q(Dout[31]), .QN(n104) );
  DF1 Dout_reg_27_ ( .D(n60), .C(Clk), .Q(Dout[27]), .QN(n26) );
  DF1 Dout_reg_26_ ( .D(n61), .C(Clk), .Q(Dout[26]), .QN(n24) );
  DF3 Dout_reg_25_ ( .D(n62), .C(Clk), .Q(Dout[25]), .QN(n22) );
  NAND23 U4 ( .A(Din[29]), .B(n317), .Q(n102) );
  NAND22 U6 ( .A(Din[24]), .B(n315), .Q(n49) );
  NAND22 U8 ( .A(Din[19]), .B(n320), .Q(n44) );
  NAND22 U10 ( .A(Dout[19]), .B(n107), .Q(n314) );
  NAND22 U12 ( .A(n314), .B(n44), .Q(n68) );
  NAND23 U14 ( .A(Din[31]), .B(n317), .Q(n105) );
  NAND23 U16 ( .A(Din[26]), .B(n316), .Q(n51) );
  NAND23 U18 ( .A(Din[30]), .B(n316), .Q(n103) );
  NAND22 U20 ( .A(Din[27]), .B(n317), .Q(n52) );
  CLKBU2 U22 ( .A(n322), .Q(n317) );
  CLKBU2 U24 ( .A(n322), .Q(n315) );
  CLKBU2 U26 ( .A(n323), .Q(n318) );
  CLKBU2 U28 ( .A(n323), .Q(n320) );
  CLKBU2 U30 ( .A(n323), .Q(n319) );
  CLKBU2 U32 ( .A(n322), .Q(n316) );
  CLKBU2 U34 ( .A(n19), .Q(n324) );
  INV3 U36 ( .A(n107), .Q(n321) );
  CLKBU2 U38 ( .A(n19), .Q(n322) );
  CLKBU2 U39 ( .A(n19), .Q(n323) );
  NAND22 U40 ( .A(Din[8]), .B(n324), .Q(n33) );
  NAND22 U42 ( .A(Din[2]), .B(n324), .Q(n21) );
  NAND22 U44 ( .A(Din[9]), .B(n318), .Q(n34) );
  NAND22 U46 ( .A(Din[7]), .B(n324), .Q(n31) );
  NAND22 U48 ( .A(Din[16]), .B(n319), .Q(n41) );
  NAND22 U50 ( .A(Din[28]), .B(n316), .Q(n101) );
  NAND22 U52 ( .A(Din[25]), .B(n317), .Q(n50) );
  NAND22 U54 ( .A(Din[17]), .B(n320), .Q(n42) );
  NAND22 U56 ( .A(Din[20]), .B(n319), .Q(n45) );
  NAND22 U58 ( .A(Din[22]), .B(n315), .Q(n47) );
  NAND22 U60 ( .A(Din[21]), .B(n315), .Q(n46) );
  NAND22 U62 ( .A(Din[23]), .B(n315), .Q(n48) );
  NAND22 U64 ( .A(Din[18]), .B(n319), .Q(n43) );
  NAND22 U66 ( .A(Din[12]), .B(n318), .Q(n37) );
  NAND22 U67 ( .A(Din[13]), .B(n320), .Q(n38) );
  NAND22 U68 ( .A(Din[14]), .B(n319), .Q(n39) );
  NAND22 U69 ( .A(Din[15]), .B(n320), .Q(n40) );
  NAND22 U70 ( .A(Din[10]), .B(n318), .Q(n35) );
  NAND22 U71 ( .A(Din[11]), .B(n318), .Q(n36) );
  NAND22 U72 ( .A(Din[6]), .B(n324), .Q(n29) );
  NAND22 U73 ( .A(Din[5]), .B(n324), .Q(n27) );
  NAND22 U74 ( .A(Din[4]), .B(n324), .Q(n25) );
  NAND22 U75 ( .A(Din[3]), .B(n324), .Q(n23) );
  NOR21 U76 ( .A(n325), .B(Reset), .Q(n19) );
  INV3 U77 ( .A(Load), .Q(n325) );
  NAND22 U78 ( .A(Din[0]), .B(n316), .Q(n106) );
  NAND22 U79 ( .A(Din[1]), .B(n324), .Q(n17) );
  NOR20 U80 ( .A(Load), .B(Reset), .Q(n107) );
endmodule


module adder_38_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n92, n97, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n418, n419, n421,
         n422, n428, n496, n569, n570, n574, n716, n717, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861;

  OAI212 U33 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U59 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n790), .C(n121), .Q(n119) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U159 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U175 ( .A(n798), .B(n790), .C(n792), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U189 ( .A(n176), .B(n790), .C(n177), .Q(n175) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  AOI212 U393 ( .A(n250), .B(n259), .C(n251), .Q(n249) );
  OAI212 U424 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U357 ( .A(n82), .B(n790), .C(n83), .Q(n81) );
  OAI212 U401 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U412 ( .A(n260), .B(n266), .C(n261), .Q(n259) );
  OAI212 U421 ( .A(n129), .B(n790), .C(n130), .Q(n128) );
  OAI212 U435 ( .A(n140), .B(n790), .C(n141), .Q(n139) );
  OAI212 U444 ( .A(n158), .B(n790), .C(n159), .Q(n157) );
  OAI212 U392 ( .A(n245), .B(n241), .C(n242), .Q(n574) );
  OAI212 U449 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U452 ( .A(n194), .B(n804), .C(n195), .Q(n191) );
  OAI212 U645 ( .A(n274), .B(n824), .C(n275), .Q(n273) );
  OAI212 U355 ( .A(n800), .B(n790), .C(n92), .Q(n90) );
  OAI212 U370 ( .A(n73), .B(n790), .C(n74), .Q(n72) );
  OAI212 U375 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  NOR24 U379 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR24 U404 ( .A(n185), .B(n194), .Q(n183) );
  XNR22 U416 ( .A(n12), .B(n90), .Q(SUM[26]) );
  AOI212 U417 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR24 U436 ( .A(B[3]), .B(A[3]), .Q(n271) );
  XNR22 U441 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U443 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U451 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U453 ( .A(n17), .B(n139), .Q(SUM[21]) );
  AOI212 U454 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  XNR22 U460 ( .A(n18), .B(n146), .Q(SUM[20]) );
  AOI212 U541 ( .A(n179), .B(n247), .C(n180), .Q(n178) );
  NOR24 U362 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR24 U366 ( .A(B[5]), .B(A[5]), .Q(n260) );
  OAI212 U380 ( .A(n158), .B(n790), .C(n159), .Q(n421) );
  OAI212 U384 ( .A(n64), .B(n790), .C(n65), .Q(n63) );
  OAI212 U385 ( .A(n801), .B(n790), .C(n795), .Q(n108) );
  OAI212 U418 ( .A(n790), .B(n102), .C(n103), .Q(n101) );
  OAI212 U456 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NOR24 U531 ( .A(B[11]), .B(A[11]), .Q(n223) );
  OAI212 U540 ( .A(n281), .B(n278), .C(n279), .Q(n496) );
  NOR24 U618 ( .A(B[9]), .B(A[9]), .Q(n241) );
  XOR22 U480 ( .A(n22), .B(n790), .Q(SUM[16]) );
  NOR24 U358 ( .A(B[10]), .B(A[10]), .Q(n230) );
  OAI212 U365 ( .A(n854), .B(n5), .C(n855), .Q(n56) );
  OAI212 U368 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  NOR24 U409 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR24 U414 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR24 U446 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR24 U448 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR24 U458 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR24 U461 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR24 U465 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR24 U466 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND23 U349 ( .A(n171), .B(n153), .Q(n151) );
  NAND22 U350 ( .A(n111), .B(n845), .Q(n102) );
  NAND24 U351 ( .A(n418), .B(n419), .Q(SUM[19]) );
  OAI211 U352 ( .A(n53), .B(n790), .C(n54), .Q(n52) );
  NOR22 U353 ( .A(n61), .B(n70), .Q(n59) );
  NOR24 U354 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND26 U356 ( .A(n825), .B(n819), .Q(n428) );
  XNR22 U359 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NOR22 U360 ( .A(B[20]), .B(A[20]), .Q(n144) );
  XNR22 U361 ( .A(n23), .B(n187), .Q(SUM[15]) );
  OAI211 U363 ( .A(n188), .B(n818), .C(n189), .Q(n187) );
  INV2 U364 ( .A(n204), .Q(n804) );
  AOI211 U367 ( .A(n789), .B(n845), .C(n848), .Q(n103) );
  AOI211 U369 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NOR22 U371 ( .A(n117), .B(n126), .Q(n115) );
  XNR22 U372 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XNR22 U373 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR22 U374 ( .A(n29), .B(n243), .Q(SUM[9]) );
  XNR22 U376 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U377 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND21 U378 ( .A(n111), .B(n84), .Q(n82) );
  CLKIN6 U381 ( .A(n112), .Q(n788) );
  INV10 U382 ( .A(n788), .Q(n789) );
  XNR22 U383 ( .A(n20), .B(n164), .Q(SUM[18]) );
  INV2 U386 ( .A(n135), .Q(n838) );
  NAND21 U387 ( .A(n799), .B(n135), .Q(n129) );
  NOR22 U388 ( .A(n137), .B(n144), .Q(n135) );
  NOR21 U389 ( .A(n88), .B(n846), .Q(n84) );
  NOR23 U390 ( .A(n113), .B(n151), .Q(n111) );
  NOR22 U391 ( .A(B[27]), .B(A[27]), .Q(n79) );
  AOI211 U394 ( .A(n794), .B(n122), .C(n123), .Q(n121) );
  NAND22 U395 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND24 U396 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND22 U397 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NOR23 U398 ( .A(n181), .B(n219), .Q(n179) );
  XOR21 U399 ( .A(n32), .B(n257), .Q(SUM[6]) );
  XNR21 U400 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NOR23 U402 ( .A(n79), .B(n88), .Q(n77) );
  NOR23 U403 ( .A(n252), .B(n255), .Q(n250) );
  INV3 U405 ( .A(n59), .Q(n854) );
  NAND22 U406 ( .A(n135), .B(n115), .Q(n113) );
  NOR22 U407 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR22 U408 ( .A(n260), .B(n265), .Q(n258) );
  NOR22 U410 ( .A(B[12]), .B(A[12]), .Q(n212) );
  AOI211 U411 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND22 U413 ( .A(n203), .B(n183), .Q(n181) );
  NOR22 U415 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR21 U419 ( .A(n801), .B(n846), .Q(n422) );
  NOR21 U420 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR22 U422 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR22 U423 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR23 U425 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U426 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NOR22 U427 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NAND22 U428 ( .A(n421), .B(n19), .Q(n418) );
  XOR21 U429 ( .A(n33), .B(n262), .Q(SUM[5]) );
  XOR21 U430 ( .A(n30), .B(n818), .Q(SUM[8]) );
  XNR21 U431 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XNR21 U432 ( .A(n27), .B(n225), .Q(SUM[11]) );
  AOI211 U433 ( .A(n794), .B(n842), .C(n843), .Q(n141) );
  OAI211 U434 ( .A(n88), .B(n849), .C(n89), .Q(n85) );
  NAND28 U437 ( .A(n428), .B(n249), .Q(n247) );
  NAND24 U438 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND24 U439 ( .A(n716), .B(n717), .Q(SUM[17]) );
  INV6 U440 ( .A(n268), .Q(n825) );
  OAI211 U442 ( .A(n219), .B(n818), .C(n220), .Q(n214) );
  OAI210 U445 ( .A(n42), .B(n790), .C(n43), .Q(n41) );
  OAI210 U447 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  NOR21 U450 ( .A(n46), .B(n6), .Q(n44) );
  CLKIN6 U455 ( .A(n175), .Q(n791) );
  AOI211 U457 ( .A(n574), .B(n812), .C(n813), .Q(n227) );
  NAND20 U459 ( .A(n239), .B(n812), .Q(n226) );
  INV1 U462 ( .A(n230), .Q(n812) );
  NOR23 U463 ( .A(B[26]), .B(A[26]), .Q(n88) );
  XNR21 U464 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND21 U467 ( .A(A[21]), .B(B[21]), .Q(n138) );
  INV3 U468 ( .A(n219), .Q(n811) );
  NAND21 U469 ( .A(n811), .B(n807), .Q(n208) );
  NAND22 U470 ( .A(n811), .B(n203), .Q(n197) );
  NAND22 U471 ( .A(n811), .B(n190), .Q(n188) );
  AOI211 U472 ( .A(n809), .B(n807), .C(n808), .Q(n209) );
  AOI211 U473 ( .A(n809), .B(n190), .C(n191), .Q(n189) );
  INV3 U474 ( .A(n220), .Q(n809) );
  OAI212 U475 ( .A(n151), .B(n790), .C(n152), .Q(n146) );
  AOI211 U476 ( .A(n825), .B(n258), .C(n259), .Q(n257) );
  INV15 U477 ( .A(n247), .Q(n818) );
  OAI212 U478 ( .A(n244), .B(n818), .C(n245), .Q(n243) );
  OAI212 U479 ( .A(n208), .B(n818), .C(n209), .Q(n207) );
  OAI212 U481 ( .A(n226), .B(n818), .C(n227), .Q(n225) );
  OAI212 U482 ( .A(n197), .B(n818), .C(n198), .Q(n196) );
  OAI212 U483 ( .A(n815), .B(n818), .C(n816), .Q(n232) );
  NOR23 U484 ( .A(n271), .B(n274), .Q(n269) );
  OAI211 U485 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  NAND24 U486 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND22 U487 ( .A(A[22]), .B(B[22]), .Q(n127) );
  INV1 U488 ( .A(n152), .Q(n794) );
  NAND21 U489 ( .A(n799), .B(n842), .Q(n140) );
  CLKIN1 U490 ( .A(n162), .Q(n832) );
  NOR21 U491 ( .A(n173), .B(n176), .Q(n171) );
  INV1 U492 ( .A(n151), .Q(n799) );
  INV0 U493 ( .A(n244), .Q(n814) );
  INV0 U494 ( .A(n79), .Q(n856) );
  NAND20 U495 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND21 U496 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NAND21 U497 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND21 U498 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND21 U499 ( .A(n111), .B(n66), .Q(n64) );
  NAND20 U500 ( .A(n807), .B(n213), .Q(n26) );
  NOR22 U501 ( .A(n99), .B(n106), .Q(n97) );
  NOR22 U502 ( .A(n241), .B(n244), .Q(n239) );
  NOR22 U503 ( .A(n155), .B(n162), .Q(n153) );
  NAND23 U504 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR21 U505 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND24 U506 ( .A(A[4]), .B(B[4]), .Q(n266) );
  INV1 U507 ( .A(n6), .Q(n847) );
  INV2 U508 ( .A(n5), .Q(n850) );
  INV3 U509 ( .A(n157), .Q(n793) );
  INV0 U510 ( .A(n70), .Q(n857) );
  NOR22 U511 ( .A(n223), .B(n230), .Q(n221) );
  CLKIN0 U512 ( .A(n212), .Q(n807) );
  INV0 U513 ( .A(n265), .Q(n822) );
  AOI210 U514 ( .A(n60), .B(n860), .C(n861), .Q(n47) );
  INV0 U515 ( .A(n176), .Q(n797) );
  XOR20 U516 ( .A(n281), .B(n37), .Q(SUM[1]) );
  XOR20 U517 ( .A(n36), .B(n824), .Q(SUM[2]) );
  INV0 U518 ( .A(n274), .Q(n841) );
  XNR20 U519 ( .A(n34), .B(n825), .Q(SUM[4]) );
  INV0 U520 ( .A(n255), .Q(n820) );
  NAND20 U521 ( .A(n820), .B(n256), .Q(n32) );
  INV0 U522 ( .A(n239), .Q(n815) );
  NAND20 U523 ( .A(n812), .B(n231), .Q(n28) );
  NAND20 U524 ( .A(n821), .B(n261), .Q(n33) );
  AOI210 U525 ( .A(n825), .B(n822), .C(n823), .Q(n262) );
  NAND20 U526 ( .A(n803), .B(n195), .Q(n24) );
  INV0 U527 ( .A(n99), .Q(n858) );
  NAND20 U528 ( .A(n858), .B(n100), .Q(n13) );
  NAND20 U529 ( .A(n856), .B(n80), .Q(n11) );
  NAND20 U530 ( .A(n59), .B(n860), .Q(n46) );
  CLKIN0 U532 ( .A(n231), .Q(n813) );
  CLKIN0 U533 ( .A(n144), .Q(n842) );
  OAI210 U534 ( .A(n126), .B(n839), .C(n127), .Q(n123) );
  NAND21 U535 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NOR22 U536 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND21 U537 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND21 U538 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND21 U539 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND21 U542 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND21 U543 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND22 U544 ( .A(A[24]), .B(B[24]), .Q(n107) );
  INV2 U545 ( .A(n38), .Q(SUM[0]) );
  INV3 U546 ( .A(n111), .Q(n801) );
  NAND22 U547 ( .A(n111), .B(n847), .Q(n73) );
  INV3 U548 ( .A(n52), .Q(n796) );
  NAND20 U549 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U550 ( .A(n422), .Q(n800) );
  NAND20 U551 ( .A(n111), .B(n55), .Q(n53) );
  AOI210 U552 ( .A(n789), .B(n55), .C(n56), .Q(n54) );
  NOR21 U553 ( .A(n854), .B(n6), .Q(n55) );
  NAND22 U554 ( .A(n97), .B(n77), .Q(n6) );
  INV3 U555 ( .A(n60), .Q(n855) );
  NAND22 U556 ( .A(n239), .B(n221), .Q(n219) );
  AOI210 U557 ( .A(n794), .B(n135), .C(n136), .Q(n130) );
  NAND22 U558 ( .A(n830), .B(n793), .Q(n419) );
  NAND22 U559 ( .A(n569), .B(n570), .Q(SUM[30]) );
  NAND22 U560 ( .A(n8), .B(n52), .Q(n569) );
  NAND22 U561 ( .A(n859), .B(n796), .Q(n570) );
  INV3 U562 ( .A(n8), .Q(n859) );
  INV3 U563 ( .A(n248), .Q(n819) );
  NAND22 U564 ( .A(n258), .B(n250), .Q(n248) );
  NAND24 U565 ( .A(n834), .B(n791), .Q(n717) );
  INV3 U566 ( .A(n21), .Q(n834) );
  NAND22 U567 ( .A(n171), .B(n832), .Q(n158) );
  NAND22 U568 ( .A(n122), .B(n799), .Q(n120) );
  INV3 U569 ( .A(n97), .Q(n846) );
  INV0 U570 ( .A(n172), .Q(n792) );
  INV0 U571 ( .A(n574), .Q(n816) );
  INV3 U572 ( .A(n19), .Q(n830) );
  NAND22 U573 ( .A(n829), .B(n242), .Q(n29) );
  INV0 U574 ( .A(n241), .Q(n829) );
  XNR21 U575 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U576 ( .A(n844), .B(n272), .Q(n35) );
  INV0 U577 ( .A(n271), .Q(n844) );
  NAND22 U578 ( .A(n810), .B(n224), .Q(n27) );
  INV0 U579 ( .A(n223), .Q(n810) );
  INV0 U580 ( .A(n194), .Q(n803) );
  NOR23 U581 ( .A(n205), .B(n212), .Q(n203) );
  NAND22 U582 ( .A(n826), .B(n279), .Q(n37) );
  INV0 U583 ( .A(n278), .Q(n826) );
  NAND22 U584 ( .A(n797), .B(n177), .Q(n22) );
  NAND20 U585 ( .A(n814), .B(n245), .Q(n30) );
  INV0 U586 ( .A(n260), .Q(n821) );
  NAND22 U587 ( .A(n841), .B(n275), .Q(n36) );
  INV0 U588 ( .A(n98), .Q(n849) );
  NAND22 U589 ( .A(n817), .B(n253), .Q(n31) );
  INV0 U590 ( .A(n252), .Q(n817) );
  XNR21 U591 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NAND22 U592 ( .A(n857), .B(n71), .Q(n10) );
  NAND22 U593 ( .A(n837), .B(n138), .Q(n17) );
  INV3 U594 ( .A(n137), .Q(n837) );
  NAND22 U595 ( .A(n853), .B(n62), .Q(n9) );
  INV3 U596 ( .A(n61), .Q(n853) );
  NAND22 U597 ( .A(n805), .B(n206), .Q(n25) );
  INV0 U598 ( .A(n205), .Q(n805) );
  NAND22 U599 ( .A(n802), .B(n186), .Q(n23) );
  INV0 U600 ( .A(n185), .Q(n802) );
  NAND22 U601 ( .A(n822), .B(n266), .Q(n34) );
  NAND22 U602 ( .A(n845), .B(n107), .Q(n14) );
  NAND22 U603 ( .A(n836), .B(n118), .Q(n15) );
  INV0 U604 ( .A(n117), .Q(n836) );
  NAND22 U605 ( .A(n832), .B(n163), .Q(n20) );
  INV0 U606 ( .A(n171), .Q(n798) );
  NAND22 U607 ( .A(n840), .B(n127), .Q(n16) );
  INV0 U608 ( .A(n126), .Q(n840) );
  NAND22 U609 ( .A(n851), .B(n89), .Q(n12) );
  INV3 U610 ( .A(n88), .Q(n851) );
  NAND22 U611 ( .A(n842), .B(n145), .Q(n18) );
  AOI210 U612 ( .A(n172), .B(n832), .C(n833), .Q(n159) );
  INV3 U613 ( .A(n163), .Q(n833) );
  NOR21 U614 ( .A(n194), .B(n806), .Q(n190) );
  INV0 U615 ( .A(n203), .Q(n806) );
  NOR21 U616 ( .A(n70), .B(n6), .Q(n66) );
  NOR21 U617 ( .A(n126), .B(n838), .Q(n122) );
  INV3 U619 ( .A(n107), .Q(n848) );
  AOI210 U620 ( .A(n789), .B(n44), .C(n45), .Q(n43) );
  INV3 U621 ( .A(n51), .Q(n861) );
  INV0 U622 ( .A(n136), .Q(n839) );
  INV3 U623 ( .A(n145), .Q(n843) );
  INV3 U624 ( .A(n213), .Q(n808) );
  NAND22 U625 ( .A(n835), .B(n174), .Q(n21) );
  INV0 U626 ( .A(n173), .Q(n835) );
  INV3 U627 ( .A(n106), .Q(n845) );
  INV3 U628 ( .A(n496), .Q(n824) );
  NAND22 U629 ( .A(n831), .B(n156), .Q(n19) );
  INV0 U630 ( .A(n155), .Q(n831) );
  INV3 U631 ( .A(n266), .Q(n823) );
  NAND22 U632 ( .A(n860), .B(n51), .Q(n8) );
  XNR21 U633 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U634 ( .A(n852), .B(n40), .Q(n7) );
  NAND22 U635 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND24 U636 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND24 U637 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND21 U638 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND21 U639 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND22 U640 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND22 U641 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND22 U642 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND22 U643 ( .A(B[5]), .B(A[5]), .Q(n261) );
  NAND22 U644 ( .A(B[3]), .B(A[3]), .Q(n272) );
  NAND20 U646 ( .A(n828), .B(n281), .Q(n38) );
  INV3 U647 ( .A(n280), .Q(n828) );
  NOR20 U648 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U649 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U650 ( .A(n50), .Q(n860) );
  NOR21 U651 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U652 ( .A(n39), .Q(n852) );
  NOR21 U653 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U654 ( .A(n175), .B(n21), .Q(n716) );
  AOI210 U655 ( .A(n809), .B(n203), .C(n204), .Q(n198) );
  AOI210 U656 ( .A(n789), .B(n97), .C(n98), .Q(n92) );
  AOI210 U657 ( .A(n789), .B(n84), .C(n85), .Q(n83) );
  INV0 U658 ( .A(n789), .Q(n795) );
  AOI210 U659 ( .A(n789), .B(n66), .C(n67), .Q(n65) );
  AOI210 U660 ( .A(n789), .B(n847), .C(n850), .Q(n74) );
  BUF15 U661 ( .A(n178), .Q(n790) );
endmodule


module adder_38 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_38_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_37_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n39, n40, n41, n42, n43, n44, n45, n48,
         n49, n50, n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82,
         n87, n88, n89, n91, n94, n95, n96, n97, n103, n104, n105, n106, n107,
         n108, n109, n112, n113, n114, n117, n118, n123, n124, n125, n126,
         n127, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n142, n144, n145, n150, n151, n152, n155, n156, n159, n160,
         n161, n164, n165, n167, n168, n169, n170, n171, n174, n175, n176,
         n177, n178, n183, n184, n185, n186, n187, n194, n195, n196, n199,
         n200, n201, n202, n203, n204, n205, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n220, n221, n222, n223, n228,
         n229, n230, n233, n234, n236, n237, n238, n239, n240, n241, n242,
         n243, n245, n246, n247, n248, n251, n252, n254, n255, n390, n393,
         n401, n409, n416, n422, n493, n494, n495, n496, n570, n571, n573,
         n648, n727, n728, n729, n732, n734, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n882, n883, n884, n885, n886, n887, n888;

  OAI212 U32 ( .A(n55), .B(n59), .C(n56), .Q(n54) );
  OAI212 U46 ( .A(n63), .B(n571), .C(n734), .Q(n62) );
  OAI212 U163 ( .A(n150), .B(n156), .C(n151), .Q(n145) );
  OAI212 U192 ( .A(n187), .B(n170), .C(n171), .Q(n169) );
  AOI212 U220 ( .A(n200), .B(n876), .C(n875), .Q(n187) );
  OAI212 U271 ( .A(n234), .B(n228), .C(n229), .Q(n223) );
  OAI212 U288 ( .A(n243), .B(n239), .C(n240), .Q(n238) );
  OAI212 U294 ( .A(n242), .B(n883), .C(n243), .Q(n241) );
  OAI212 U301 ( .A(n246), .B(n248), .C(n247), .Q(n245) );
  OAI212 U334 ( .A(n205), .B(n201), .C(n202), .Q(n200) );
  OAI212 U345 ( .A(n869), .B(n860), .C(n866), .Q(n196) );
  OAI212 U351 ( .A(n177), .B(n860), .C(n178), .Q(n176) );
  OAI212 U424 ( .A(n843), .B(n70), .C(n71), .Q(n69) );
  OAI212 U466 ( .A(n834), .B(n843), .C(n91), .Q(n89) );
  OAI212 U467 ( .A(n842), .B(n843), .C(n840), .Q(n114) );
  OAI212 U468 ( .A(n108), .B(n843), .C(n109), .Q(n107) );
  OAI212 U469 ( .A(n79), .B(n843), .C(n80), .Q(n78) );
  OAI212 U386 ( .A(n843), .B(n126), .C(n127), .Q(n125) );
  OAI212 U436 ( .A(n217), .B(n859), .C(n220), .Q(n216) );
  OAI212 U382 ( .A(n130), .B(n167), .C(n131), .Q(n409) );
  OAI212 U449 ( .A(n130), .B(n167), .C(n131), .Q(n129) );
  OAI212 U408 ( .A(n186), .B(n860), .C(n187), .Q(n185) );
  OAI212 U409 ( .A(n220), .B(n212), .C(n213), .Q(n211) );
  OAI212 U442 ( .A(n142), .B(n134), .C(n135), .Q(n133) );
  AOI212 U354 ( .A(n409), .B(n61), .C(n62), .Q(n1) );
  OAI212 U464 ( .A(n648), .B(n63), .C(n734), .Q(n495) );
  OAI212 U473 ( .A(n45), .B(n41), .C(n42), .Q(n40) );
  OAI212 U355 ( .A(n187), .B(n170), .C(n171), .Q(n729) );
  NAND26 U323 ( .A(n117), .B(n103), .Q(n97) );
  NOR24 U324 ( .A(n134), .B(n139), .Q(n132) );
  NAND21 U325 ( .A(B[6]), .B(A[6]), .Q(n229) );
  NOR23 U326 ( .A(A[6]), .B(B[6]), .Q(n228) );
  NAND22 U327 ( .A(B[10]), .B(A[10]), .Q(n202) );
  NOR21 U328 ( .A(A[29]), .B(B[29]), .Q(n48) );
  OAI212 U329 ( .A(n1), .B(n818), .C(n819), .Q(n36) );
  CLKIN6 U330 ( .A(n159), .Q(n854) );
  NAND26 U331 ( .A(n871), .B(n878), .Q(n170) );
  INV6 U332 ( .A(n183), .Q(n878) );
  NAND23 U333 ( .A(n810), .B(n811), .Q(n812) );
  NOR23 U335 ( .A(A[18]), .B(B[18]), .Q(n134) );
  INV3 U336 ( .A(n39), .Q(n818) );
  INV3 U337 ( .A(n390), .Q(n861) );
  NOR22 U338 ( .A(n186), .B(n170), .Q(n168) );
  NOR22 U339 ( .A(A[21]), .B(B[21]), .Q(n112) );
  NAND22 U340 ( .A(n53), .B(n822), .Q(n44) );
  NOR23 U341 ( .A(A[22]), .B(B[22]), .Q(n105) );
  INV3 U342 ( .A(n113), .Q(n839) );
  NAND22 U343 ( .A(n732), .B(n124), .Q(n493) );
  INV3 U344 ( .A(n81), .Q(n832) );
  INV3 U346 ( .A(n416), .Q(n835) );
  NOR22 U347 ( .A(A[28]), .B(B[28]), .Q(n55) );
  NOR23 U348 ( .A(A[30]), .B(B[30]), .Q(n41) );
  NAND23 U349 ( .A(n422), .B(n68), .Q(n66) );
  NOR23 U350 ( .A(n55), .B(n58), .Q(n53) );
  INV3 U352 ( .A(n48), .Q(n822) );
  NOR21 U353 ( .A(n217), .B(n212), .Q(n210) );
  NOR22 U356 ( .A(A[9]), .B(B[9]), .Q(n204) );
  NAND23 U357 ( .A(n199), .B(n876), .Q(n186) );
  INV3 U358 ( .A(n144), .Q(n848) );
  NOR22 U359 ( .A(A[19]), .B(B[19]), .Q(n126) );
  NAND22 U360 ( .A(A[21]), .B(B[21]), .Q(n113) );
  INV3 U361 ( .A(n41), .Q(n817) );
  NAND22 U362 ( .A(B[27]), .B(A[27]), .Q(n59) );
  AOI211 U363 ( .A(n880), .B(n222), .C(n223), .Q(n221) );
  NAND22 U364 ( .A(B[9]), .B(A[9]), .Q(n205) );
  NAND23 U365 ( .A(B[19]), .B(A[19]), .Q(n127) );
  INV3 U366 ( .A(n2), .Q(n814) );
  XOR21 U367 ( .A(n15), .B(n136), .Q(SUM[18]) );
  NAND24 U368 ( .A(A[20]), .B(n813), .Q(n124) );
  INV3 U369 ( .A(n82), .Q(n831) );
  INV6 U370 ( .A(n87), .Q(n811) );
  INV2 U371 ( .A(n160), .Q(n855) );
  NAND22 U372 ( .A(n854), .B(n160), .Q(n18) );
  NAND22 U373 ( .A(B[15]), .B(A[15]), .Q(n160) );
  OAI210 U374 ( .A(n390), .B(n848), .C(n846), .Q(n393) );
  CLKIN3 U375 ( .A(n201), .Q(n868) );
  NOR21 U376 ( .A(n204), .B(n201), .Q(n199) );
  NOR23 U377 ( .A(A[10]), .B(B[10]), .Q(n201) );
  NAND24 U378 ( .A(n812), .B(n88), .Q(n82) );
  INV6 U379 ( .A(n95), .Q(n810) );
  NAND24 U380 ( .A(n570), .B(n124), .Q(n118) );
  INV2 U381 ( .A(n97), .Q(n837) );
  INV2 U383 ( .A(n494), .Q(n834) );
  NAND21 U384 ( .A(n129), .B(n837), .Q(n573) );
  NAND24 U385 ( .A(n836), .B(n839), .Q(n401) );
  NAND24 U387 ( .A(n850), .B(n841), .Q(n570) );
  INV6 U388 ( .A(n127), .Q(n850) );
  CLKIN3 U389 ( .A(n74), .Q(n830) );
  CLKIN1 U390 ( .A(n134), .Q(n849) );
  CLKIN0 U391 ( .A(n117), .Q(n842) );
  NAND20 U392 ( .A(n117), .B(n838), .Q(n108) );
  NAND23 U393 ( .A(B[23]), .B(A[23]), .Q(n95) );
  NOR24 U394 ( .A(A[23]), .B(B[23]), .Q(n94) );
  INV0 U395 ( .A(n126), .Q(n851) );
  NOR24 U396 ( .A(A[26]), .B(B[26]), .Q(n67) );
  NAND22 U397 ( .A(B[12]), .B(A[12]), .Q(n184) );
  INV2 U398 ( .A(n94), .Q(n833) );
  INV3 U399 ( .A(n207), .Q(n860) );
  AOI211 U400 ( .A(n207), .B(n168), .C(n729), .Q(n390) );
  OAI212 U401 ( .A(n208), .B(n236), .C(n209), .Q(n207) );
  NOR22 U402 ( .A(A[12]), .B(B[12]), .Q(n183) );
  NOR24 U403 ( .A(B[20]), .B(A[20]), .Q(n123) );
  BUF12 U404 ( .A(B[20]), .Q(n813) );
  NOR22 U405 ( .A(n123), .B(n126), .Q(n117) );
  INV3 U406 ( .A(n49), .Q(n820) );
  NAND20 U407 ( .A(n822), .B(n49), .Q(n4) );
  NAND22 U410 ( .A(B[28]), .B(A[28]), .Q(n56) );
  NOR23 U411 ( .A(n41), .B(n44), .Q(n39) );
  NAND22 U412 ( .A(B[30]), .B(A[30]), .Q(n42) );
  CLKIN6 U413 ( .A(n67), .Q(n828) );
  NAND21 U414 ( .A(n837), .B(n81), .Q(n79) );
  NOR20 U415 ( .A(n97), .B(n94), .Q(n494) );
  NAND22 U416 ( .A(B[29]), .B(A[29]), .Q(n49) );
  NAND28 U417 ( .A(n401), .B(n106), .Q(n104) );
  NOR22 U418 ( .A(A[7]), .B(B[7]), .Q(n217) );
  NOR24 U419 ( .A(n63), .B(n97), .Q(n61) );
  NAND22 U420 ( .A(A[22]), .B(B[22]), .Q(n106) );
  INV1 U421 ( .A(n112), .Q(n838) );
  NOR23 U422 ( .A(n74), .B(n67), .Q(n65) );
  CLKIN6 U423 ( .A(n105), .Q(n836) );
  INV1 U425 ( .A(n145), .Q(n846) );
  NAND21 U426 ( .A(B[26]), .B(A[26]), .Q(n68) );
  NAND21 U427 ( .A(n823), .B(n56), .Q(n5) );
  NOR22 U428 ( .A(B[15]), .B(A[15]), .Q(n159) );
  NOR22 U429 ( .A(n150), .B(n155), .Q(n144) );
  NAND21 U430 ( .A(n573), .B(n416), .Q(n96) );
  NOR22 U431 ( .A(A[13]), .B(B[13]), .Q(n174) );
  XOR22 U432 ( .A(n814), .B(n36), .Q(SUM[31]) );
  NOR23 U433 ( .A(B[25]), .B(A[25]), .Q(n74) );
  NAND22 U434 ( .A(B[25]), .B(A[25]), .Q(n77) );
  NAND21 U435 ( .A(n838), .B(n113), .Q(n12) );
  CLKIN3 U437 ( .A(n53), .Q(n825) );
  CLKIN6 U438 ( .A(n123), .Q(n841) );
  AOI212 U439 ( .A(n871), .B(n877), .C(n872), .Q(n171) );
  INV3 U440 ( .A(n175), .Q(n872) );
  NOR24 U441 ( .A(n112), .B(n105), .Q(n103) );
  INV0 U443 ( .A(n139), .Q(n844) );
  NOR20 U444 ( .A(n139), .B(n848), .Q(n137) );
  NOR23 U445 ( .A(A[17]), .B(B[17]), .Q(n139) );
  OAI211 U446 ( .A(n204), .B(n860), .C(n205), .Q(n203) );
  NAND22 U447 ( .A(A[17]), .B(B[17]), .Q(n142) );
  NOR24 U448 ( .A(A[24]), .B(B[24]), .Q(n87) );
  NAND21 U450 ( .A(A[18]), .B(B[18]), .Q(n135) );
  AOI212 U451 ( .A(n118), .B(n103), .C(n104), .Q(n648) );
  CLKIN2 U452 ( .A(n50), .Q(n824) );
  OAI212 U453 ( .A(n825), .B(n496), .C(n826), .Q(n50) );
  AOI211 U454 ( .A(n835), .B(n833), .C(n810), .Q(n91) );
  AOI211 U455 ( .A(n835), .B(n72), .C(n73), .Q(n71) );
  INV0 U456 ( .A(n55), .Q(n823) );
  NAND24 U457 ( .A(n132), .B(n144), .Q(n130) );
  XOR20 U458 ( .A(n6), .B(n1), .Q(SUM[27]) );
  NAND21 U459 ( .A(B[13]), .B(A[13]), .Q(n175) );
  NOR24 U460 ( .A(n815), .B(A[16]), .Q(n150) );
  AOI212 U461 ( .A(n118), .B(n103), .C(n104), .Q(n571) );
  AOI212 U462 ( .A(n245), .B(n237), .C(n238), .Q(n236) );
  AOI212 U463 ( .A(n854), .B(n856), .C(n855), .Q(n156) );
  NAND21 U465 ( .A(n830), .B(n77), .Q(n8) );
  OAI210 U470 ( .A(n74), .B(n831), .C(n77), .Q(n73) );
  CLKIN3 U471 ( .A(n77), .Q(n829) );
  NOR24 U472 ( .A(n94), .B(n87), .Q(n81) );
  BUF6 U474 ( .A(B[16]), .Q(n815) );
  AOI212 U475 ( .A(n132), .B(n145), .C(n133), .Q(n131) );
  AOI211 U476 ( .A(n861), .B(n857), .C(n856), .Q(n161) );
  NAND26 U477 ( .A(n65), .B(n81), .Q(n63) );
  AOI212 U478 ( .A(n822), .B(n54), .C(n820), .Q(n45) );
  OAI210 U479 ( .A(n139), .B(n846), .C(n142), .Q(n138) );
  NAND21 U480 ( .A(A[24]), .B(B[24]), .Q(n88) );
  INV2 U481 ( .A(n58), .Q(n827) );
  NOR22 U482 ( .A(B[27]), .B(A[27]), .Q(n58) );
  AOI212 U483 ( .A(n103), .B(n493), .C(n104), .Q(n416) );
  OAI211 U484 ( .A(n496), .B(n58), .C(n59), .Q(n57) );
  AOI212 U485 ( .A(n409), .B(n61), .C(n495), .Q(n496) );
  AOI211 U486 ( .A(n835), .B(n81), .C(n82), .Q(n80) );
  AOI212 U487 ( .A(n65), .B(n82), .C(n66), .Q(n734) );
  NAND21 U488 ( .A(n833), .B(n95), .Q(n10) );
  NAND21 U489 ( .A(n50), .B(n4), .Q(n727) );
  INV0 U490 ( .A(n493), .Q(n840) );
  INV2 U491 ( .A(n4), .Q(n821) );
  AOI212 U492 ( .A(n207), .B(n168), .C(n169), .Q(n167) );
  CLKIN0 U493 ( .A(n222), .Q(n863) );
  NAND21 U494 ( .A(B[7]), .B(A[7]), .Q(n220) );
  NAND21 U495 ( .A(B[11]), .B(A[11]), .Q(n195) );
  INV3 U496 ( .A(n174), .Q(n871) );
  NAND22 U497 ( .A(B[5]), .B(A[5]), .Q(n234) );
  NAND21 U498 ( .A(n817), .B(n42), .Q(n3) );
  XNR20 U499 ( .A(n19), .B(n861), .Q(SUM[14]) );
  CLKIN0 U500 ( .A(n54), .Q(n826) );
  INV0 U501 ( .A(n155), .Q(n853) );
  INV0 U502 ( .A(n156), .Q(n852) );
  INV0 U503 ( .A(n199), .Q(n869) );
  INV0 U504 ( .A(n236), .Q(n880) );
  INV0 U505 ( .A(n223), .Q(n859) );
  NAND21 U506 ( .A(n837), .B(n72), .Q(n70) );
  AOI211 U507 ( .A(n137), .B(n861), .C(n138), .Q(n136) );
  NOR20 U508 ( .A(n217), .B(n863), .Q(n215) );
  INV0 U509 ( .A(n186), .Q(n870) );
  NAND20 U510 ( .A(n878), .B(n870), .Q(n177) );
  AOI210 U511 ( .A(n867), .B(n878), .C(n877), .Q(n178) );
  INV0 U512 ( .A(n217), .Q(n864) );
  INV0 U513 ( .A(n233), .Q(n862) );
  INV0 U514 ( .A(n150), .Q(n847) );
  INV0 U515 ( .A(n228), .Q(n865) );
  INV0 U516 ( .A(n204), .Q(n873) );
  NAND20 U517 ( .A(n879), .B(n240), .Q(n29) );
  INV0 U518 ( .A(n212), .Q(n874) );
  NAND20 U519 ( .A(B[8]), .B(A[8]), .Q(n213) );
  NOR20 U520 ( .A(A[4]), .B(B[4]), .Q(n239) );
  NAND21 U521 ( .A(B[31]), .B(A[31]), .Q(n35) );
  INV2 U522 ( .A(n34), .Q(n816) );
  NAND20 U523 ( .A(n874), .B(n213), .Q(n25) );
  INV6 U524 ( .A(n129), .Q(n843) );
  INV3 U525 ( .A(n393), .Q(n845) );
  INV0 U526 ( .A(n200), .Q(n866) );
  AOI211 U527 ( .A(n861), .B(n853), .C(n852), .Q(n152) );
  INV0 U528 ( .A(n187), .Q(n867) );
  INV3 U529 ( .A(n245), .Q(n883) );
  INV3 U530 ( .A(n195), .Q(n875) );
  NAND22 U531 ( .A(n222), .B(n210), .Q(n208) );
  AOI211 U532 ( .A(n223), .B(n210), .C(n211), .Q(n209) );
  NOR21 U533 ( .A(n242), .B(n239), .Q(n237) );
  NOR21 U534 ( .A(n228), .B(n233), .Q(n222) );
  INV3 U535 ( .A(n40), .Q(n819) );
  AOI211 U536 ( .A(n880), .B(n215), .C(n216), .Q(n214) );
  AOI211 U537 ( .A(n880), .B(n862), .C(n858), .Q(n230) );
  INV3 U538 ( .A(n234), .Q(n858) );
  NAND22 U539 ( .A(n857), .B(n854), .Q(n155) );
  NAND22 U540 ( .A(n850), .B(n841), .Q(n732) );
  NAND22 U541 ( .A(n829), .B(n828), .Q(n422) );
  INV3 U542 ( .A(n242), .Q(n887) );
  INV3 U543 ( .A(n184), .Q(n877) );
  INV3 U544 ( .A(n165), .Q(n856) );
  INV3 U545 ( .A(n239), .Q(n879) );
  INV3 U546 ( .A(n246), .Q(n888) );
  AOI211 U547 ( .A(n885), .B(n884), .C(n886), .Q(n248) );
  INV3 U548 ( .A(n252), .Q(n886) );
  NOR21 U549 ( .A(A[3]), .B(B[3]), .Q(n242) );
  NOR21 U550 ( .A(A[8]), .B(B[8]), .Q(n212) );
  NOR21 U551 ( .A(A[5]), .B(B[5]), .Q(n233) );
  NAND22 U552 ( .A(B[14]), .B(A[14]), .Q(n165) );
  NAND22 U553 ( .A(n815), .B(A[16]), .Q(n151) );
  NAND22 U554 ( .A(B[4]), .B(A[4]), .Q(n240) );
  INV3 U555 ( .A(n194), .Q(n876) );
  NOR21 U556 ( .A(A[11]), .B(B[11]), .Q(n194) );
  INV3 U557 ( .A(n164), .Q(n857) );
  NOR21 U558 ( .A(A[14]), .B(B[14]), .Q(n164) );
  NOR21 U559 ( .A(A[2]), .B(B[2]), .Q(n246) );
  INV3 U560 ( .A(n251), .Q(n885) );
  NOR21 U561 ( .A(A[1]), .B(B[1]), .Q(n251) );
  NAND22 U562 ( .A(B[1]), .B(A[1]), .Q(n252) );
  NAND22 U563 ( .A(B[3]), .B(A[3]), .Q(n243) );
  NAND22 U564 ( .A(B[2]), .B(A[2]), .Q(n247) );
  INV3 U565 ( .A(n255), .Q(n884) );
  NOR21 U566 ( .A(A[31]), .B(B[31]), .Q(n34) );
  INV3 U567 ( .A(n254), .Q(n882) );
  NOR21 U568 ( .A(A[0]), .B(B[0]), .Q(n254) );
  NAND22 U569 ( .A(B[0]), .B(A[0]), .Q(n255) );
  XNR21 U570 ( .A(n11), .B(n107), .Q(SUM[22]) );
  NAND20 U571 ( .A(n836), .B(n106), .Q(n11) );
  XNR21 U572 ( .A(n8), .B(n78), .Q(SUM[25]) );
  XNR21 U573 ( .A(n13), .B(n125), .Q(SUM[20]) );
  NAND20 U574 ( .A(n124), .B(n841), .Q(n13) );
  XNR21 U575 ( .A(n7), .B(n69), .Q(SUM[26]) );
  NAND20 U576 ( .A(n68), .B(n828), .Q(n7) );
  XNR21 U577 ( .A(n5), .B(n57), .Q(SUM[28]) );
  NAND22 U578 ( .A(n816), .B(n35), .Q(n2) );
  XNR21 U579 ( .A(n10), .B(n96), .Q(SUM[23]) );
  XOR20 U580 ( .A(n14), .B(n843), .Q(SUM[19]) );
  NAND20 U581 ( .A(n851), .B(n127), .Q(n14) );
  XOR21 U582 ( .A(n16), .B(n845), .Q(SUM[17]) );
  NAND20 U583 ( .A(n844), .B(n142), .Q(n16) );
  XOR21 U584 ( .A(n17), .B(n152), .Q(SUM[16]) );
  NAND20 U585 ( .A(n847), .B(n151), .Q(n17) );
  XNR21 U586 ( .A(n20), .B(n176), .Q(SUM[13]) );
  NAND20 U587 ( .A(n871), .B(n175), .Q(n20) );
  XNR21 U588 ( .A(n23), .B(n203), .Q(SUM[10]) );
  NAND20 U589 ( .A(n868), .B(n202), .Q(n23) );
  XNR21 U590 ( .A(n22), .B(n196), .Q(SUM[11]) );
  NAND20 U591 ( .A(n876), .B(n195), .Q(n22) );
  NAND20 U592 ( .A(n857), .B(n165), .Q(n19) );
  XOR21 U593 ( .A(n26), .B(n221), .Q(SUM[7]) );
  NAND20 U594 ( .A(n864), .B(n220), .Q(n26) );
  XOR21 U595 ( .A(n25), .B(n214), .Q(SUM[8]) );
  XNR21 U596 ( .A(n3), .B(n43), .Q(SUM[30]) );
  XNR21 U597 ( .A(n12), .B(n114), .Q(SUM[21]) );
  XNR21 U598 ( .A(n9), .B(n89), .Q(SUM[24]) );
  NAND20 U599 ( .A(n811), .B(n88), .Q(n9) );
  NAND20 U600 ( .A(n827), .B(n59), .Q(n6) );
  NAND20 U601 ( .A(n849), .B(n135), .Q(n15) );
  XOR21 U602 ( .A(n18), .B(n161), .Q(SUM[15]) );
  XNR21 U603 ( .A(n21), .B(n185), .Q(SUM[12]) );
  NAND20 U604 ( .A(n878), .B(n184), .Q(n21) );
  XOR21 U605 ( .A(n30), .B(n883), .Q(SUM[3]) );
  NAND22 U606 ( .A(n887), .B(n243), .Q(n30) );
  XOR21 U607 ( .A(n27), .B(n230), .Q(SUM[6]) );
  NAND20 U608 ( .A(n865), .B(n229), .Q(n27) );
  XOR21 U609 ( .A(n24), .B(n860), .Q(SUM[9]) );
  NAND20 U610 ( .A(n873), .B(n205), .Q(n24) );
  NAND22 U611 ( .A(n727), .B(n728), .Q(SUM[29]) );
  NAND22 U612 ( .A(n824), .B(n821), .Q(n728) );
  XNR21 U613 ( .A(n884), .B(n32), .Q(SUM[1]) );
  NAND22 U614 ( .A(n885), .B(n252), .Q(n32) );
  XOR21 U615 ( .A(n31), .B(n248), .Q(SUM[2]) );
  NAND22 U616 ( .A(n888), .B(n247), .Q(n31) );
  XNR21 U617 ( .A(n29), .B(n241), .Q(SUM[4]) );
  XNR21 U618 ( .A(n28), .B(n880), .Q(SUM[5]) );
  NAND20 U619 ( .A(n862), .B(n234), .Q(n28) );
  INV3 U620 ( .A(n33), .Q(SUM[0]) );
  NAND22 U621 ( .A(n882), .B(n255), .Q(n33) );
  NOR21 U622 ( .A(n74), .B(n832), .Q(n72) );
  OAI211 U623 ( .A(n1), .B(n44), .C(n45), .Q(n43) );
  AOI210 U624 ( .A(n493), .B(n838), .C(n839), .Q(n109) );
endmodule


module adder_37 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_37_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_36_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n420, n556, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n817, n818, n819, n820, n821, n822;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U101 ( .A(n776), .B(n759), .C(n774), .Q(n108) );
  OAI212 U115 ( .A(n120), .B(n759), .C(n121), .Q(n119) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U175 ( .A(n785), .B(n759), .C(n782), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U233 ( .A(n208), .B(n789), .C(n209), .Q(n207) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U257 ( .A(n226), .B(n789), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n793), .B(n789), .C(n795), .Q(n232) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n818), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U420 ( .A(n140), .B(n759), .C(n141), .Q(n139) );
  OAI212 U422 ( .A(n158), .B(n759), .C(n159), .Q(n157) );
  OAI212 U423 ( .A(n102), .B(n759), .C(n103), .Q(n101) );
  OAI212 U354 ( .A(n73), .B(n759), .C(n74), .Q(n72) );
  OAI212 U461 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U407 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U395 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U485 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U435 ( .A(n197), .B(n789), .C(n198), .Q(n196) );
  OAI212 U478 ( .A(n213), .B(n205), .C(n556), .Q(n420) );
  OAI212 U367 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U413 ( .A(n42), .B(n759), .C(n43), .Q(n41) );
  OAI212 U408 ( .A(n91), .B(n759), .C(n92), .Q(n90) );
  OAI212 U370 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U421 ( .A(n82), .B(n759), .C(n83), .Q(n81) );
  OAI212 U433 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U441 ( .A(n219), .B(n789), .C(n220), .Q(n214) );
  OAI212 U458 ( .A(n126), .B(n781), .C(n127), .Q(n123) );
  XNR22 U349 ( .A(n28), .B(n232), .Q(SUM[10]) );
  AOI212 U350 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  OAI211 U351 ( .A(n205), .B(n213), .C(n556), .Q(n204) );
  NOR23 U352 ( .A(n185), .B(n194), .Q(n183) );
  NOR24 U353 ( .A(B[14]), .B(A[14]), .Q(n194) );
  OAI210 U355 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  NAND21 U356 ( .A(A[21]), .B(B[21]), .Q(n138) );
  XNR22 U357 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XNR22 U358 ( .A(n29), .B(n243), .Q(SUM[9]) );
  OAI212 U359 ( .A(n244), .B(n789), .C(n245), .Q(n243) );
  XNR22 U360 ( .A(n17), .B(n139), .Q(SUM[21]) );
  AOI210 U361 ( .A(n783), .B(n135), .C(n136), .Q(n130) );
  INV2 U362 ( .A(n152), .Q(n783) );
  NOR23 U363 ( .A(n113), .B(n151), .Q(n111) );
  NAND24 U364 ( .A(n171), .B(n153), .Q(n151) );
  XNR22 U365 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NOR21 U366 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U368 ( .A(n88), .B(n772), .Q(n84) );
  INV3 U369 ( .A(n97), .Q(n772) );
  NOR21 U371 ( .A(n173), .B(n176), .Q(n171) );
  NOR23 U372 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR21 U373 ( .A(B[28]), .B(A[28]), .Q(n70) );
  INV1 U374 ( .A(n212), .Q(n803) );
  INV3 U375 ( .A(n244), .Q(n811) );
  NOR22 U376 ( .A(n79), .B(n88), .Q(n77) );
  NOR22 U377 ( .A(n117), .B(n126), .Q(n115) );
  NOR22 U378 ( .A(n137), .B(n144), .Q(n135) );
  NOR23 U379 ( .A(n155), .B(n162), .Q(n153) );
  NAND22 U380 ( .A(n203), .B(n183), .Q(n181) );
  INV3 U381 ( .A(n98), .Q(n773) );
  NOR21 U382 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR23 U383 ( .A(n205), .B(n212), .Q(n203) );
  NAND22 U384 ( .A(A[16]), .B(B[16]), .Q(n177) );
  XNR21 U385 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XNR21 U386 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR21 U387 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NOR24 U388 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR22 U389 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND20 U390 ( .A(n556), .B(n815), .Q(n25) );
  NOR23 U391 ( .A(B[11]), .B(A[11]), .Q(n223) );
  OAI211 U392 ( .A(n194), .B(n806), .C(n195), .Q(n191) );
  NAND22 U393 ( .A(n786), .B(n135), .Q(n129) );
  NOR23 U394 ( .A(B[22]), .B(A[22]), .Q(n126) );
  OAI211 U396 ( .A(n64), .B(n759), .C(n65), .Q(n63) );
  NOR24 U397 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR23 U398 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NAND21 U399 ( .A(B[13]), .B(A[13]), .Q(n556) );
  NOR21 U400 ( .A(n765), .B(n6), .Q(n55) );
  NOR24 U401 ( .A(B[15]), .B(A[15]), .Q(n185) );
  XOR22 U402 ( .A(n22), .B(n759), .Q(SUM[16]) );
  NOR23 U403 ( .A(B[12]), .B(A[12]), .Q(n212) );
  XNR22 U404 ( .A(n23), .B(n187), .Q(SUM[15]) );
  OAI211 U405 ( .A(n188), .B(n789), .C(n189), .Q(n187) );
  OAI210 U406 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  CLKIN3 U409 ( .A(n5), .Q(n768) );
  OAI211 U410 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  NAND21 U411 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND21 U412 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NOR21 U414 ( .A(B[7]), .B(A[7]), .Q(n252) );
  XNR22 U415 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND22 U416 ( .A(n111), .B(n84), .Q(n82) );
  OAI212 U417 ( .A(n151), .B(n759), .C(n152), .Q(n146) );
  AOI211 U418 ( .A(n758), .B(n66), .C(n67), .Q(n65) );
  NAND22 U419 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NAND22 U424 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NOR22 U425 ( .A(B[27]), .B(A[27]), .Q(n79) );
  OAI212 U426 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  XNR22 U427 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NOR24 U428 ( .A(B[13]), .B(A[13]), .Q(n205) );
  AOI211 U429 ( .A(n783), .B(n778), .C(n780), .Q(n141) );
  INV0 U430 ( .A(n144), .Q(n778) );
  XNR22 U431 ( .A(n15), .B(n119), .Q(SUM[23]) );
  AOI211 U432 ( .A(n758), .B(n769), .C(n768), .Q(n74) );
  BUF12 U434 ( .A(n112), .Q(n758) );
  NOR22 U436 ( .A(B[18]), .B(A[18]), .Q(n162) );
  XNR22 U437 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U438 ( .A(n12), .B(n90), .Q(SUM[26]) );
  AOI211 U439 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NAND21 U440 ( .A(A[19]), .B(B[19]), .Q(n156) );
  XNR22 U442 ( .A(n18), .B(n146), .Q(SUM[20]) );
  INV3 U443 ( .A(n162), .Q(n798) );
  XNR22 U444 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND21 U445 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NOR20 U446 ( .A(n252), .B(n255), .Q(n250) );
  OAI211 U447 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U448 ( .A(n129), .B(n759), .C(n130), .Q(n128) );
  OAI212 U449 ( .A(n88), .B(n773), .C(n89), .Q(n85) );
  NAND21 U450 ( .A(A[26]), .B(B[26]), .Q(n89) );
  XNR22 U451 ( .A(n9), .B(n63), .Q(SUM[29]) );
  CLKIN2 U452 ( .A(n203), .Q(n804) );
  XNR22 U453 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U454 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND21 U455 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NOR20 U456 ( .A(n241), .B(n244), .Q(n239) );
  NAND21 U457 ( .A(A[23]), .B(B[23]), .Q(n118) );
  XNR22 U459 ( .A(n21), .B(n175), .Q(SUM[17]) );
  OAI211 U460 ( .A(n176), .B(n759), .C(n177), .Q(n175) );
  OAI212 U462 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  INV1 U463 ( .A(n107), .Q(n800) );
  NAND22 U464 ( .A(A[20]), .B(B[20]), .Q(n145) );
  INV1 U465 ( .A(n137), .Q(n797) );
  NOR21 U466 ( .A(B[29]), .B(A[29]), .Q(n61) );
  OAI210 U467 ( .A(n53), .B(n759), .C(n54), .Q(n52) );
  NAND21 U468 ( .A(n810), .B(n186), .Q(n23) );
  NAND21 U469 ( .A(A[15]), .B(B[15]), .Q(n186) );
  CLKIN3 U470 ( .A(n117), .Q(n775) );
  OAI211 U471 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  BUF15 U472 ( .A(n178), .Q(n759) );
  NOR22 U473 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR22 U474 ( .A(n99), .B(n106), .Q(n97) );
  INV2 U475 ( .A(n99), .Q(n771) );
  AOI211 U476 ( .A(n758), .B(n97), .C(n98), .Q(n92) );
  NAND22 U477 ( .A(n111), .B(n97), .Q(n91) );
  INV2 U479 ( .A(n205), .Q(n815) );
  NOR22 U480 ( .A(B[16]), .B(A[16]), .Q(n176) );
  INV0 U481 ( .A(n185), .Q(n810) );
  INV2 U482 ( .A(n106), .Q(n801) );
  INV2 U483 ( .A(n151), .Q(n786) );
  NAND21 U484 ( .A(n788), .B(n261), .Q(n33) );
  NAND20 U486 ( .A(n814), .B(n224), .Q(n27) );
  INV3 U487 ( .A(n6), .Q(n769) );
  INV3 U488 ( .A(n220), .Q(n796) );
  NOR23 U489 ( .A(n181), .B(n219), .Q(n179) );
  NAND22 U490 ( .A(n792), .B(n242), .Q(n29) );
  INV2 U491 ( .A(n241), .Q(n792) );
  NAND22 U492 ( .A(n807), .B(n253), .Q(n31) );
  INV2 U493 ( .A(n252), .Q(n807) );
  NAND20 U494 ( .A(n798), .B(n163), .Q(n20) );
  NAND20 U495 ( .A(n813), .B(n174), .Q(n21) );
  CLKIN1 U496 ( .A(n758), .Q(n774) );
  NAND20 U497 ( .A(n801), .B(n107), .Q(n14) );
  NAND22 U498 ( .A(n811), .B(n245), .Q(n30) );
  NAND22 U499 ( .A(n812), .B(n256), .Q(n32) );
  INV2 U500 ( .A(n255), .Q(n812) );
  INV3 U501 ( .A(n265), .Q(n791) );
  NAND22 U502 ( .A(n111), .B(n801), .Q(n102) );
  CLKIN3 U503 ( .A(n60), .Q(n764) );
  OAI210 U504 ( .A(n765), .B(n5), .C(n764), .Q(n56) );
  AOI210 U505 ( .A(n796), .B(n203), .C(n420), .Q(n198) );
  NAND20 U506 ( .A(n794), .B(n203), .Q(n197) );
  NAND20 U507 ( .A(n794), .B(n190), .Q(n188) );
  AOI211 U508 ( .A(n758), .B(n801), .C(n800), .Q(n103) );
  INV0 U509 ( .A(n136), .Q(n781) );
  INV0 U510 ( .A(n155), .Q(n802) );
  INV0 U511 ( .A(n126), .Q(n777) );
  NAND20 U512 ( .A(n777), .B(n127), .Q(n16) );
  AOI210 U513 ( .A(n60), .B(n762), .C(n761), .Q(n47) );
  NAND20 U514 ( .A(n784), .B(n177), .Q(n22) );
  AOI211 U515 ( .A(n796), .B(n803), .C(n805), .Q(n209) );
  INV0 U516 ( .A(n213), .Q(n805) );
  INV0 U517 ( .A(n194), .Q(n787) );
  NAND20 U518 ( .A(n767), .B(n80), .Q(n11) );
  NAND20 U519 ( .A(n239), .B(n808), .Q(n226) );
  CLKIN3 U520 ( .A(n239), .Q(n793) );
  NOR21 U521 ( .A(n61), .B(n70), .Q(n59) );
  INV0 U522 ( .A(n70), .Q(n766) );
  NAND21 U523 ( .A(n766), .B(n71), .Q(n10) );
  INV0 U524 ( .A(n173), .Q(n813) );
  CLKIN0 U525 ( .A(n171), .Q(n785) );
  NAND20 U526 ( .A(n803), .B(n213), .Q(n26) );
  NOR20 U527 ( .A(n260), .B(n265), .Q(n258) );
  NOR20 U528 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NOR20 U529 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR21 U530 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND20 U531 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND20 U532 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND20 U533 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U534 ( .A(n111), .B(n769), .Q(n73) );
  INV3 U535 ( .A(n111), .Q(n776) );
  NAND20 U536 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U537 ( .A(n219), .Q(n794) );
  NAND22 U538 ( .A(n97), .B(n77), .Q(n6) );
  NOR20 U539 ( .A(n46), .B(n6), .Q(n44) );
  NAND20 U540 ( .A(n111), .B(n66), .Q(n64) );
  NAND22 U541 ( .A(n135), .B(n115), .Q(n113) );
  INV3 U542 ( .A(n59), .Q(n765) );
  NAND22 U543 ( .A(n786), .B(n122), .Q(n120) );
  NAND21 U544 ( .A(n786), .B(n778), .Q(n140) );
  NAND22 U545 ( .A(n171), .B(n798), .Q(n158) );
  INV0 U546 ( .A(n172), .Q(n782) );
  AOI211 U547 ( .A(n819), .B(n258), .C(n259), .Q(n257) );
  NAND22 U548 ( .A(n239), .B(n221), .Q(n219) );
  INV3 U549 ( .A(n247), .Q(n789) );
  INV3 U550 ( .A(n268), .Q(n819) );
  INV3 U551 ( .A(n277), .Q(n818) );
  NAND22 U552 ( .A(n794), .B(n803), .Q(n208) );
  INV3 U553 ( .A(n240), .Q(n795) );
  XOR21 U554 ( .A(n30), .B(n789), .Q(SUM[8]) );
  XOR21 U555 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U556 ( .A(n819), .B(n791), .C(n790), .Q(n262) );
  INV3 U557 ( .A(n266), .Q(n790) );
  INV3 U558 ( .A(n176), .Q(n784) );
  NAND22 U559 ( .A(n762), .B(n51), .Q(n8) );
  NAND20 U560 ( .A(n111), .B(n55), .Q(n53) );
  NAND22 U561 ( .A(n763), .B(n62), .Q(n9) );
  INV3 U562 ( .A(n61), .Q(n763) );
  NAND20 U563 ( .A(n787), .B(n195), .Q(n24) );
  NAND22 U564 ( .A(n808), .B(n231), .Q(n28) );
  XNR21 U565 ( .A(n34), .B(n819), .Q(SUM[4]) );
  NAND22 U566 ( .A(n791), .B(n266), .Q(n34) );
  XNR21 U567 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U568 ( .A(n771), .B(n100), .Q(n13) );
  XNR21 U569 ( .A(n11), .B(n81), .Q(SUM[27]) );
  INV0 U570 ( .A(n79), .Q(n767) );
  NAND22 U571 ( .A(n778), .B(n145), .Q(n18) );
  INV3 U572 ( .A(n51), .Q(n761) );
  NOR21 U573 ( .A(n70), .B(n6), .Q(n66) );
  NAND20 U574 ( .A(n797), .B(n138), .Q(n17) );
  NAND22 U575 ( .A(n775), .B(n118), .Q(n15) );
  NOR21 U576 ( .A(n126), .B(n779), .Q(n122) );
  INV0 U577 ( .A(n135), .Q(n779) );
  NAND20 U578 ( .A(n802), .B(n156), .Q(n19) );
  NAND22 U579 ( .A(n770), .B(n89), .Q(n12) );
  INV3 U580 ( .A(n88), .Q(n770) );
  NOR21 U581 ( .A(n194), .B(n804), .Q(n190) );
  AOI211 U582 ( .A(n796), .B(n190), .C(n191), .Q(n189) );
  INV3 U583 ( .A(n420), .Q(n806) );
  AOI211 U584 ( .A(n783), .B(n122), .C(n123), .Q(n121) );
  AOI210 U585 ( .A(n172), .B(n798), .C(n799), .Q(n159) );
  INV3 U586 ( .A(n163), .Q(n799) );
  INV3 U587 ( .A(n145), .Q(n780) );
  NAND21 U588 ( .A(n59), .B(n762), .Q(n46) );
  INV3 U589 ( .A(n230), .Q(n808) );
  INV3 U590 ( .A(n223), .Q(n814) );
  INV3 U591 ( .A(n260), .Q(n788) );
  XOR21 U592 ( .A(n32), .B(n257), .Q(SUM[6]) );
  XOR21 U593 ( .A(n36), .B(n818), .Q(SUM[2]) );
  NAND22 U594 ( .A(n821), .B(n275), .Q(n36) );
  INV3 U595 ( .A(n274), .Q(n821) );
  XOR21 U596 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U597 ( .A(n820), .B(n279), .Q(n37) );
  INV3 U598 ( .A(n278), .Q(n820) );
  XNR21 U599 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U600 ( .A(n822), .B(n272), .Q(n35) );
  INV3 U601 ( .A(n271), .Q(n822) );
  AOI211 U602 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U603 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U604 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U605 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U606 ( .A(n223), .B(n230), .Q(n221) );
  AOI210 U607 ( .A(n240), .B(n808), .C(n809), .Q(n227) );
  INV3 U608 ( .A(n231), .Q(n809) );
  NAND22 U609 ( .A(B[12]), .B(A[12]), .Q(n213) );
  XNR21 U610 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U611 ( .A(n760), .B(n40), .Q(n7) );
  NAND21 U612 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND20 U613 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NOR22 U614 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR21 U615 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV3 U616 ( .A(n50), .Q(n762) );
  NAND20 U617 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV3 U618 ( .A(n39), .Q(n760) );
  NOR20 U619 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND20 U620 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND20 U621 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND20 U622 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND20 U623 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND20 U624 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV3 U625 ( .A(n38), .Q(SUM[0]) );
  NAND22 U626 ( .A(n817), .B(n281), .Q(n38) );
  INV3 U627 ( .A(n280), .Q(n817) );
  NOR20 U628 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NOR20 U629 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR20 U630 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND20 U631 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U632 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NOR20 U633 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND20 U634 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U635 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U636 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND20 U637 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NOR20 U638 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NOR21 U639 ( .A(B[24]), .B(A[24]), .Q(n106) );
  AOI210 U640 ( .A(n758), .B(n44), .C(n45), .Q(n43) );
  AOI210 U641 ( .A(n758), .B(n55), .C(n56), .Q(n54) );
  AOI210 U642 ( .A(n758), .B(n84), .C(n85), .Q(n83) );
endmodule


module adder_36 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_36_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_35_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n232, n239, n240, n241, n242, n243, n244, n245, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n265, n266, n268, n269, n270, n271, n272, n273,
         n274, n275, n277, n278, n279, n280, n281, n429, n431, n498, n641,
         n642, n714, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U91 ( .A(n102), .B(n799), .C(n103), .Q(n101) );
  OAI212 U101 ( .A(n431), .B(n799), .C(n839), .Q(n108) );
  OAI212 U127 ( .A(n129), .B(n799), .C(n130), .Q(n128) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n799), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U175 ( .A(n850), .B(n799), .C(n852), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U233 ( .A(n208), .B(n804), .C(n209), .Q(n207) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U257 ( .A(n226), .B(n804), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n816), .B(n804), .C(n818), .Q(n232) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n802), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U422 ( .A(n188), .B(n804), .C(n189), .Q(n187) );
  OAI212 U438 ( .A(n158), .B(n799), .C(n159), .Q(n157) );
  OAI212 U367 ( .A(n197), .B(n804), .C(n198), .Q(n196) );
  OAI212 U472 ( .A(n120), .B(n799), .C(n121), .Q(n119) );
  OAI212 U486 ( .A(n91), .B(n799), .C(n92), .Q(n90) );
  OAI212 U452 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U445 ( .A(n42), .B(n799), .C(n43), .Q(n41) );
  OAI212 U465 ( .A(n714), .B(n223), .C(n224), .Q(n222) );
  OAI212 U455 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U401 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U421 ( .A(n151), .B(n799), .C(n152), .Q(n146) );
  OAI212 U396 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U413 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U429 ( .A(n89), .B(n798), .C(n80), .Q(n78) );
  XNR22 U349 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND21 U350 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND22 U351 ( .A(n203), .B(n183), .Q(n181) );
  NOR23 U352 ( .A(n185), .B(n194), .Q(n183) );
  INV2 U353 ( .A(n204), .Q(n857) );
  NAND21 U354 ( .A(B[21]), .B(A[21]), .Q(n138) );
  NAND21 U355 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NOR24 U356 ( .A(A[11]), .B(B[11]), .Q(n223) );
  XNR22 U357 ( .A(n28), .B(n232), .Q(SUM[10]) );
  CLKIN6 U358 ( .A(n112), .Q(n786) );
  NAND21 U359 ( .A(A[23]), .B(B[23]), .Q(n118) );
  AOI211 U360 ( .A(n853), .B(n135), .C(n136), .Q(n130) );
  NOR24 U361 ( .A(A[13]), .B(B[13]), .Q(n205) );
  NOR23 U362 ( .A(B[12]), .B(A[12]), .Q(n212) );
  XNR22 U363 ( .A(n19), .B(n157), .Q(SUM[19]) );
  CLKIN12 U364 ( .A(n786), .Q(n787) );
  XNR22 U365 ( .A(n17), .B(n139), .Q(SUM[21]) );
  NAND21 U366 ( .A(n851), .B(n847), .Q(n140) );
  INV6 U368 ( .A(n151), .Q(n851) );
  NAND24 U369 ( .A(n842), .B(n851), .Q(n431) );
  NOR21 U370 ( .A(n194), .B(n856), .Q(n190) );
  INV1 U371 ( .A(n203), .Q(n856) );
  INV3 U372 ( .A(n108), .Q(n790) );
  XNR21 U373 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NOR22 U374 ( .A(n155), .B(n162), .Q(n153) );
  NOR22 U375 ( .A(n798), .B(n88), .Q(n77) );
  NOR22 U376 ( .A(n99), .B(n106), .Q(n97) );
  NOR22 U377 ( .A(B[18]), .B(A[18]), .Q(n162) );
  CLKIN3 U378 ( .A(n128), .Q(n794) );
  NOR22 U379 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND22 U380 ( .A(n841), .B(n84), .Q(n82) );
  XNR21 U381 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NOR23 U382 ( .A(B[15]), .B(A[15]), .Q(n185) );
  AOI211 U383 ( .A(n819), .B(n190), .C(n191), .Q(n189) );
  INV3 U384 ( .A(n247), .Q(n804) );
  NAND24 U385 ( .A(n791), .B(n792), .Q(SUM[24]) );
  NAND24 U386 ( .A(n789), .B(n790), .Q(n792) );
  XNR21 U387 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XOR21 U388 ( .A(n32), .B(n257), .Q(SUM[6]) );
  OAI211 U389 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  INV3 U390 ( .A(n137), .Q(n797) );
  NAND21 U391 ( .A(n841), .B(n55), .Q(n53) );
  INV3 U392 ( .A(n787), .Q(n839) );
  INV2 U393 ( .A(n839), .Q(n788) );
  NAND21 U394 ( .A(n797), .B(n138), .Q(n17) );
  NOR23 U395 ( .A(n137), .B(n144), .Q(n135) );
  INV2 U397 ( .A(n144), .Q(n847) );
  NAND21 U398 ( .A(n851), .B(n135), .Q(n129) );
  NAND28 U399 ( .A(n641), .B(n642), .Q(SUM[20]) );
  NAND24 U400 ( .A(n845), .B(n806), .Q(n642) );
  NOR22 U402 ( .A(n173), .B(n176), .Q(n171) );
  NOR23 U403 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR24 U404 ( .A(B[17]), .B(A[17]), .Q(n173) );
  INV0 U405 ( .A(n714), .Q(n862) );
  NAND22 U406 ( .A(n14), .B(n108), .Q(n791) );
  INV3 U407 ( .A(n14), .Q(n789) );
  NOR22 U408 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND22 U409 ( .A(n837), .B(n107), .Q(n14) );
  NOR21 U410 ( .A(B[8]), .B(A[8]), .Q(n244) );
  AOI211 U411 ( .A(n819), .B(n203), .C(n204), .Q(n198) );
  AOI212 U412 ( .A(n183), .B(n204), .C(n184), .Q(n182) );
  AOI210 U414 ( .A(n787), .B(n66), .C(n67), .Q(n65) );
  OAI211 U415 ( .A(n64), .B(n799), .C(n65), .Q(n63) );
  NAND21 U416 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NOR21 U417 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND22 U418 ( .A(n498), .B(n83), .Q(n81) );
  INV2 U419 ( .A(n136), .Q(n846) );
  OAI212 U420 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  NAND22 U423 ( .A(n832), .B(n805), .Q(n498) );
  INV1 U424 ( .A(n799), .Q(n805) );
  OAI211 U425 ( .A(n53), .B(n799), .C(n54), .Q(n52) );
  NAND22 U426 ( .A(n16), .B(n128), .Q(n795) );
  NAND24 U427 ( .A(n793), .B(n794), .Q(n796) );
  NAND28 U428 ( .A(n795), .B(n796), .Q(SUM[22]) );
  INV6 U430 ( .A(n16), .Q(n793) );
  NAND22 U431 ( .A(n843), .B(n127), .Q(n16) );
  INV2 U432 ( .A(n152), .Q(n853) );
  NAND21 U433 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NOR22 U434 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR24 U435 ( .A(A[14]), .B(B[14]), .Q(n194) );
  NOR21 U436 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND23 U437 ( .A(n135), .B(n115), .Q(n113) );
  XOR21 U439 ( .A(n22), .B(n799), .Q(SUM[16]) );
  OAI212 U440 ( .A(n176), .B(n799), .C(n177), .Q(n175) );
  OAI212 U441 ( .A(n194), .B(n857), .C(n195), .Q(n191) );
  AOI212 U442 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NOR22 U443 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR22 U444 ( .A(n117), .B(n126), .Q(n115) );
  OAI212 U446 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NAND22 U447 ( .A(A[12]), .B(B[12]), .Q(n213) );
  INV3 U448 ( .A(n82), .Q(n832) );
  NOR21 U449 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NOR20 U450 ( .A(n223), .B(n230), .Q(n221) );
  INV1 U451 ( .A(n223), .Q(n854) );
  AOI212 U453 ( .A(n787), .B(n97), .C(n98), .Q(n92) );
  NOR21 U454 ( .A(n70), .B(n6), .Q(n66) );
  XNR22 U456 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NOR20 U457 ( .A(B[2]), .B(A[2]), .Q(n274) );
  OAI212 U458 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  NAND22 U459 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND22 U460 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND21 U461 ( .A(A[24]), .B(B[24]), .Q(n107) );
  INV10 U462 ( .A(n431), .Q(n841) );
  CLKIN1 U463 ( .A(n135), .Q(n848) );
  OAI211 U464 ( .A(n73), .B(n799), .C(n74), .Q(n72) );
  INV1 U466 ( .A(n117), .Q(n840) );
  AOI210 U467 ( .A(n787), .B(n84), .C(n85), .Q(n83) );
  NOR20 U468 ( .A(B[10]), .B(A[10]), .Q(n230) );
  XNR22 U469 ( .A(n23), .B(n187), .Q(SUM[15]) );
  XNR22 U470 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NOR23 U471 ( .A(n205), .B(n212), .Q(n203) );
  NAND22 U473 ( .A(n863), .B(n714), .Q(n28) );
  NAND22 U474 ( .A(A[10]), .B(B[10]), .Q(n714) );
  XNR22 U475 ( .A(n15), .B(n119), .Q(SUM[23]) );
  XNR22 U476 ( .A(n13), .B(n101), .Q(SUM[25]) );
  OAI211 U477 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI210 U478 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  NOR20 U479 ( .A(n241), .B(n244), .Q(n239) );
  OAI210 U480 ( .A(n244), .B(n804), .C(n245), .Q(n243) );
  CLKIN2 U481 ( .A(n244), .Q(n815) );
  XNR22 U482 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NOR21 U483 ( .A(B[28]), .B(A[28]), .Q(n70) );
  XNR22 U484 ( .A(n12), .B(n90), .Q(SUM[26]) );
  BUF6 U485 ( .A(n79), .Q(n798) );
  BUF15 U487 ( .A(n178), .Q(n799) );
  NAND21 U488 ( .A(n841), .B(n830), .Q(n73) );
  NAND21 U489 ( .A(n841), .B(n66), .Q(n64) );
  XNR22 U490 ( .A(n11), .B(n81), .Q(SUM[27]) );
  INV0 U491 ( .A(n173), .Q(n849) );
  NAND21 U492 ( .A(A[20]), .B(B[20]), .Q(n145) );
  INV1 U493 ( .A(n145), .Q(n844) );
  AOI212 U494 ( .A(n787), .B(n837), .C(n838), .Q(n103) );
  AOI211 U495 ( .A(n787), .B(n830), .C(n828), .Q(n74) );
  NOR21 U496 ( .A(B[24]), .B(A[24]), .Q(n106) );
  INV2 U497 ( .A(n126), .Q(n843) );
  OAI210 U498 ( .A(n126), .B(n846), .C(n127), .Q(n123) );
  INV1 U499 ( .A(n155), .Q(n860) );
  NOR23 U500 ( .A(A[19]), .B(B[19]), .Q(n155) );
  INV2 U501 ( .A(n212), .Q(n866) );
  NOR21 U502 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NAND22 U503 ( .A(n18), .B(n146), .Q(n641) );
  CLKIN2 U504 ( .A(n97), .Q(n834) );
  NAND22 U505 ( .A(A[16]), .B(B[16]), .Q(n177) );
  CLKIN2 U506 ( .A(n18), .Q(n845) );
  INV3 U507 ( .A(n220), .Q(n819) );
  INV0 U508 ( .A(n172), .Q(n852) );
  NAND22 U509 ( .A(n827), .B(n71), .Q(n10) );
  NAND22 U510 ( .A(n97), .B(n851), .Q(n429) );
  NAND21 U511 ( .A(n835), .B(n842), .Q(n91) );
  OAI210 U512 ( .A(n826), .B(n5), .C(n825), .Q(n56) );
  NAND22 U513 ( .A(n820), .B(n242), .Q(n29) );
  INV2 U514 ( .A(n241), .Q(n820) );
  INV0 U515 ( .A(n70), .Q(n827) );
  NAND20 U516 ( .A(n831), .B(n89), .Q(n12) );
  CLKIN1 U517 ( .A(n98), .Q(n836) );
  OAI211 U518 ( .A(n88), .B(n836), .C(n89), .Q(n85) );
  NAND22 U519 ( .A(n815), .B(n245), .Q(n30) );
  INV2 U520 ( .A(n265), .Q(n810) );
  NOR20 U521 ( .A(n826), .B(n6), .Q(n55) );
  NOR22 U522 ( .A(n181), .B(n219), .Q(n179) );
  NAND22 U523 ( .A(n171), .B(n153), .Q(n151) );
  CLKIN3 U524 ( .A(n60), .Q(n825) );
  INV3 U525 ( .A(n5), .Q(n828) );
  CLKIN3 U526 ( .A(n59), .Q(n826) );
  NAND20 U527 ( .A(n817), .B(n203), .Q(n197) );
  AOI211 U528 ( .A(n819), .B(n866), .C(n867), .Q(n209) );
  INV0 U529 ( .A(n213), .Q(n867) );
  INV0 U530 ( .A(n88), .Q(n831) );
  NAND20 U531 ( .A(n866), .B(n213), .Q(n26) );
  AOI211 U532 ( .A(n240), .B(n863), .C(n862), .Q(n227) );
  CLKIN3 U533 ( .A(n239), .Q(n816) );
  AOI210 U534 ( .A(n853), .B(n847), .C(n844), .Q(n141) );
  NAND22 U535 ( .A(n812), .B(n261), .Q(n33) );
  NAND20 U536 ( .A(n847), .B(n145), .Q(n18) );
  NAND21 U537 ( .A(n59), .B(n823), .Q(n46) );
  NAND20 U538 ( .A(n858), .B(n163), .Q(n20) );
  INV0 U539 ( .A(n61), .Q(n824) );
  INV3 U540 ( .A(n230), .Q(n863) );
  INV0 U541 ( .A(n185), .Q(n865) );
  NAND20 U542 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U543 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND20 U544 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U545 ( .A(A[4]), .B(B[4]), .Q(n266) );
  INV3 U546 ( .A(n146), .Q(n806) );
  NAND20 U547 ( .A(n841), .B(n44), .Q(n42) );
  INV3 U548 ( .A(n113), .Q(n842) );
  INV3 U549 ( .A(n6), .Q(n830) );
  INV3 U550 ( .A(n219), .Q(n817) );
  NAND22 U551 ( .A(n97), .B(n77), .Q(n6) );
  NOR20 U552 ( .A(n46), .B(n6), .Q(n44) );
  NAND20 U553 ( .A(n171), .B(n858), .Q(n158) );
  NAND21 U554 ( .A(n851), .B(n122), .Q(n120) );
  NAND22 U555 ( .A(n841), .B(n837), .Q(n102) );
  CLKIN0 U556 ( .A(n171), .Q(n850) );
  INV3 U557 ( .A(n429), .Q(n835) );
  AOI211 U558 ( .A(n803), .B(n258), .C(n259), .Q(n257) );
  NAND22 U559 ( .A(n239), .B(n221), .Q(n219) );
  INV3 U560 ( .A(n268), .Q(n803) );
  INV3 U561 ( .A(n277), .Q(n802) );
  INV3 U562 ( .A(n240), .Q(n818) );
  NAND22 U563 ( .A(n239), .B(n863), .Q(n226) );
  NAND22 U564 ( .A(n817), .B(n190), .Q(n188) );
  NAND22 U565 ( .A(n817), .B(n866), .Q(n208) );
  NAND22 U566 ( .A(n864), .B(n177), .Q(n22) );
  INV0 U567 ( .A(n176), .Q(n864) );
  XOR21 U568 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U569 ( .A(n803), .B(n810), .C(n811), .Q(n262) );
  INV3 U570 ( .A(n266), .Q(n811) );
  NAND22 U571 ( .A(n813), .B(n256), .Q(n32) );
  INV2 U572 ( .A(n255), .Q(n813) );
  XOR21 U573 ( .A(n30), .B(n804), .Q(SUM[8]) );
  AOI210 U574 ( .A(n60), .B(n823), .C(n822), .Q(n47) );
  INV3 U575 ( .A(n51), .Q(n822) );
  INV3 U576 ( .A(n107), .Q(n838) );
  NAND22 U577 ( .A(n833), .B(n100), .Q(n13) );
  INV3 U578 ( .A(n99), .Q(n833) );
  NAND20 U579 ( .A(n865), .B(n186), .Q(n23) );
  NAND22 U580 ( .A(n829), .B(n80), .Q(n11) );
  INV3 U581 ( .A(n798), .Q(n829) );
  XNR21 U582 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND22 U583 ( .A(n824), .B(n62), .Q(n9) );
  NAND20 U584 ( .A(n849), .B(n174), .Q(n21) );
  XNR21 U585 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND22 U586 ( .A(n823), .B(n51), .Q(n8) );
  NAND20 U587 ( .A(n206), .B(n855), .Q(n25) );
  INV3 U588 ( .A(n205), .Q(n855) );
  XNR21 U589 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U590 ( .A(n224), .B(n854), .Q(n27) );
  XNR21 U591 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U592 ( .A(n809), .B(n272), .Q(n35) );
  INV3 U593 ( .A(n271), .Q(n809) );
  NAND22 U594 ( .A(n814), .B(n253), .Q(n31) );
  INV3 U595 ( .A(n252), .Q(n814) );
  XNR21 U596 ( .A(n34), .B(n803), .Q(SUM[4]) );
  NAND22 U597 ( .A(n810), .B(n266), .Q(n34) );
  XNR21 U598 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NOR21 U599 ( .A(n61), .B(n70), .Q(n59) );
  NAND22 U600 ( .A(n840), .B(n118), .Q(n15) );
  NOR21 U601 ( .A(n88), .B(n834), .Q(n84) );
  NAND20 U602 ( .A(n860), .B(n156), .Q(n19) );
  NOR21 U603 ( .A(n126), .B(n848), .Q(n122) );
  NAND20 U604 ( .A(n861), .B(n195), .Q(n24) );
  INV3 U605 ( .A(n194), .Q(n861) );
  AOI210 U606 ( .A(n172), .B(n858), .C(n859), .Q(n159) );
  INV3 U607 ( .A(n163), .Q(n859) );
  CLKIN3 U608 ( .A(n260), .Q(n812) );
  AOI211 U609 ( .A(n853), .B(n122), .C(n123), .Q(n121) );
  INV3 U610 ( .A(n162), .Q(n858) );
  INV3 U611 ( .A(n106), .Q(n837) );
  XOR21 U612 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U613 ( .A(n807), .B(n279), .Q(n37) );
  INV3 U614 ( .A(n278), .Q(n807) );
  XOR21 U615 ( .A(n36), .B(n802), .Q(SUM[2]) );
  NAND22 U616 ( .A(n808), .B(n275), .Q(n36) );
  INV3 U617 ( .A(n274), .Q(n808) );
  AOI211 U618 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U619 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U620 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U621 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR20 U622 ( .A(n252), .B(n255), .Q(n250) );
  NOR20 U623 ( .A(n260), .B(n265), .Q(n258) );
  XNR21 U624 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U625 ( .A(n821), .B(n40), .Q(n7) );
  NAND20 U626 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR20 U627 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NAND21 U628 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND20 U629 ( .A(A[28]), .B(B[28]), .Q(n71) );
  INV3 U630 ( .A(n50), .Q(n823) );
  NOR20 U631 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U632 ( .A(n39), .Q(n821) );
  NOR20 U633 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U634 ( .A(n38), .Q(SUM[0]) );
  NAND22 U635 ( .A(n801), .B(n281), .Q(n38) );
  INV3 U636 ( .A(n280), .Q(n801) );
  NOR20 U637 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U638 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U639 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND20 U640 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND20 U641 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U642 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U643 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND20 U644 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NOR20 U645 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NAND21 U646 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND22 U647 ( .A(B[14]), .B(A[14]), .Q(n195) );
  NAND20 U648 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NOR21 U649 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND20 U650 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NOR21 U651 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND21 U652 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NOR21 U653 ( .A(B[1]), .B(A[1]), .Q(n278) );
  OAI210 U654 ( .A(n219), .B(n804), .C(n220), .Q(n214) );
  NOR22 U655 ( .A(B[26]), .B(A[26]), .Q(n88) );
  AOI210 U656 ( .A(n788), .B(n44), .C(n45), .Q(n43) );
  AOI210 U657 ( .A(n787), .B(n55), .C(n56), .Q(n54) );
  NOR21 U658 ( .A(B[7]), .B(A[7]), .Q(n252) );
endmodule


module adder_35 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_35_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_34_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n74, n78, n79, n80, n81, n82, n83, n84, n85,
         n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103, n106,
         n107, n108, n111, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n126, n127, n128, n129, n130, n135, n136, n137,
         n138, n139, n140, n141, n144, n145, n146, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n162, n163, n164, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n194, n195, n196, n197,
         n198, n203, n204, n205, n206, n207, n208, n209, n212, n213, n214,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n230, n231,
         n232, n239, n240, n241, n242, n243, n244, n245, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n265, n266, n268, n269, n270, n271, n272, n273, n274,
         n275, n277, n278, n279, n280, n281, n422, n423, n425, n439, n507,
         n516, n592, n604, n673, n674, n756, n758, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n911, n912, n913;

  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  AOI212 U157 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n911), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U352 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U379 ( .A(n208), .B(n886), .C(n209), .Q(n207) );
  OAI212 U381 ( .A(n226), .B(n886), .C(n227), .Q(n225) );
  OAI212 U382 ( .A(n894), .B(n886), .C(n892), .Q(n232) );
  OAI212 U386 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U395 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U437 ( .A(n120), .B(n843), .C(n121), .Q(n119) );
  OAI212 U474 ( .A(n856), .B(n843), .C(n74), .Q(n72) );
  AOI212 U542 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI212 U483 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U503 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  AOI212 U665 ( .A(n874), .B(n866), .C(n864), .Q(n604) );
  OAI212 U384 ( .A(n244), .B(n886), .C(n245), .Q(n243) );
  OAI212 U487 ( .A(n843), .B(n102), .C(n103), .Q(n101) );
  OAI212 U502 ( .A(n155), .B(n163), .C(n156), .Q(n154) );
  OAI212 U518 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U427 ( .A(n188), .B(n886), .C(n189), .Q(n187) );
  OAI212 U465 ( .A(n197), .B(n886), .C(n198), .Q(n196) );
  OAI212 U484 ( .A(n176), .B(n843), .C(n177), .Q(n175) );
  OAI212 U485 ( .A(n158), .B(n843), .C(n159), .Q(n157) );
  OAI212 U494 ( .A(n861), .B(n88), .C(n89), .Q(n85) );
  NAND20 U349 ( .A(n891), .B(n203), .Q(n197) );
  NAND22 U350 ( .A(B[12]), .B(A[12]), .Q(n213) );
  NOR24 U351 ( .A(n162), .B(n155), .Q(n153) );
  CLKIN6 U353 ( .A(n152), .Q(n874) );
  NAND22 U354 ( .A(B[13]), .B(A[13]), .Q(n206) );
  NOR23 U355 ( .A(n46), .B(n6), .Q(n44) );
  NAND23 U356 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND28 U357 ( .A(n203), .B(n183), .Q(n181) );
  CLKIN3 U358 ( .A(n60), .Q(n847) );
  AOI212 U359 ( .A(n60), .B(n845), .C(n846), .Q(n47) );
  NOR24 U360 ( .A(n223), .B(n230), .Q(n221) );
  NOR22 U361 ( .A(A[11]), .B(B[11]), .Q(n223) );
  AOI211 U362 ( .A(n863), .B(n44), .C(n45), .Q(n43) );
  INV3 U363 ( .A(n113), .Q(n866) );
  NAND28 U364 ( .A(n135), .B(n115), .Q(n113) );
  NOR24 U365 ( .A(n117), .B(n126), .Q(n115) );
  NAND21 U366 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NOR22 U367 ( .A(B[14]), .B(A[14]), .Q(n194) );
  XNR22 U368 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NOR24 U369 ( .A(A[22]), .B(B[22]), .Q(n126) );
  NAND23 U370 ( .A(n171), .B(n153), .Q(n151) );
  AOI212 U371 ( .A(n863), .B(n97), .C(n674), .Q(n92) );
  CLKIN2 U372 ( .A(n863), .Q(n841) );
  NAND21 U373 ( .A(n876), .B(n881), .Q(n140) );
  NOR24 U374 ( .A(n185), .B(n194), .Q(n183) );
  INV1 U375 ( .A(n106), .Q(n858) );
  NAND22 U376 ( .A(n111), .B(n834), .Q(n835) );
  INV3 U377 ( .A(n14), .Q(n830) );
  NOR22 U378 ( .A(A[24]), .B(B[24]), .Q(n106) );
  NOR22 U380 ( .A(n867), .B(n6), .Q(n758) );
  INV3 U383 ( .A(n843), .Q(n884) );
  INV3 U385 ( .A(n874), .Q(n836) );
  NOR23 U387 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR23 U388 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR22 U389 ( .A(n173), .B(n176), .Q(n171) );
  NOR23 U390 ( .A(A[15]), .B(B[15]), .Q(n185) );
  NOR22 U391 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U392 ( .A(A[28]), .B(B[28]), .Q(n71) );
  INV3 U393 ( .A(n70), .Q(n851) );
  NAND23 U394 ( .A(n239), .B(n221), .Q(n219) );
  NAND22 U396 ( .A(A[16]), .B(B[16]), .Q(n177) );
  XNR21 U397 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR21 U398 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR21 U399 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND22 U400 ( .A(n111), .B(n858), .Q(n102) );
  NAND22 U401 ( .A(A[17]), .B(B[17]), .Q(n174) );
  INV2 U402 ( .A(n889), .Q(n829) );
  INV3 U403 ( .A(n220), .Q(n889) );
  CLKIN1 U404 ( .A(n205), .Q(n898) );
  AOI211 U405 ( .A(n837), .B(n135), .C(n842), .Q(n130) );
  INV3 U406 ( .A(n162), .Q(n875) );
  XNR21 U407 ( .A(n20), .B(n164), .Q(SUM[18]) );
  CLKIN6 U408 ( .A(n117), .Q(n865) );
  OAI211 U409 ( .A(n129), .B(n843), .C(n130), .Q(n128) );
  INV2 U410 ( .A(n151), .Q(n876) );
  INV0 U411 ( .A(n185), .Q(n885) );
  CLKIN3 U412 ( .A(n111), .Q(n867) );
  NAND21 U413 ( .A(n14), .B(n108), .Q(n832) );
  NAND22 U414 ( .A(n830), .B(n831), .Q(n833) );
  NAND22 U415 ( .A(n832), .B(n833), .Q(SUM[24]) );
  CLKIN6 U416 ( .A(n108), .Q(n831) );
  NAND26 U417 ( .A(n835), .B(n841), .Q(n108) );
  INV3 U418 ( .A(n843), .Q(n834) );
  NAND24 U419 ( .A(n868), .B(n865), .Q(n439) );
  NAND23 U420 ( .A(n439), .B(n118), .Q(n116) );
  OAI210 U421 ( .A(n219), .B(n886), .C(n829), .Q(n214) );
  NAND24 U422 ( .A(n673), .B(n54), .Q(n52) );
  AOI212 U423 ( .A(n863), .B(n55), .C(n56), .Q(n54) );
  NOR23 U424 ( .A(n850), .B(n6), .Q(n55) );
  NAND21 U425 ( .A(n111), .B(n44), .Q(n42) );
  NAND21 U426 ( .A(n111), .B(n66), .Q(n64) );
  NAND21 U428 ( .A(n111), .B(n55), .Q(n53) );
  INV3 U429 ( .A(n758), .Q(n856) );
  INV8 U430 ( .A(n604), .Q(n863) );
  INV0 U431 ( .A(n223), .Q(n903) );
  INV3 U432 ( .A(n842), .Q(n870) );
  OAI211 U433 ( .A(n137), .B(n145), .C(n138), .Q(n842) );
  AOI211 U434 ( .A(n837), .B(n122), .C(n123), .Q(n121) );
  NOR21 U435 ( .A(n126), .B(n872), .Q(n122) );
  OAI211 U436 ( .A(n516), .B(n850), .C(n847), .Q(n56) );
  OAI212 U438 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  INV1 U439 ( .A(n203), .Q(n899) );
  NOR24 U440 ( .A(A[13]), .B(B[13]), .Q(n205) );
  INV3 U441 ( .A(n836), .Q(n837) );
  NAND22 U442 ( .A(n838), .B(n839), .Q(n840) );
  NAND23 U443 ( .A(n840), .B(n92), .Q(n90) );
  INV3 U444 ( .A(n91), .Q(n838) );
  INV2 U445 ( .A(n843), .Q(n839) );
  NAND24 U446 ( .A(n849), .B(n884), .Q(n673) );
  AOI212 U447 ( .A(n863), .B(n858), .C(n860), .Q(n103) );
  OAI212 U448 ( .A(n140), .B(n843), .C(n141), .Q(n139) );
  AOI210 U449 ( .A(n889), .B(n203), .C(n425), .Q(n198) );
  AOI212 U450 ( .A(n863), .B(n84), .C(n85), .Q(n83) );
  CLKIN4 U451 ( .A(n114), .Q(n864) );
  OAI212 U452 ( .A(n137), .B(n145), .C(n138), .Q(n136) );
  CLKIN3 U453 ( .A(n194), .Q(n902) );
  OAI210 U454 ( .A(n194), .B(n897), .C(n195), .Q(n191) );
  NOR20 U455 ( .A(n194), .B(n899), .Q(n190) );
  AOI212 U456 ( .A(n863), .B(n66), .C(n67), .Q(n65) );
  NAND21 U457 ( .A(B[15]), .B(A[15]), .Q(n186) );
  OAI211 U458 ( .A(n151), .B(n843), .C(n836), .Q(n146) );
  NOR23 U459 ( .A(n219), .B(n181), .Q(n179) );
  CLKIN6 U460 ( .A(n5), .Q(n853) );
  NAND21 U461 ( .A(n111), .B(n84), .Q(n82) );
  AOI212 U462 ( .A(n863), .B(n855), .C(n853), .Q(n74) );
  INV1 U463 ( .A(n6), .Q(n855) );
  XNR22 U464 ( .A(n7), .B(n41), .Q(SUM[31]) );
  CLKIN0 U466 ( .A(n163), .Q(n873) );
  NAND21 U467 ( .A(B[11]), .B(A[11]), .Q(n224) );
  NAND22 U468 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND21 U469 ( .A(n845), .B(n51), .Q(n8) );
  NAND21 U470 ( .A(A[30]), .B(B[30]), .Q(n51) );
  XNR22 U471 ( .A(n12), .B(n90), .Q(SUM[26]) );
  INV2 U472 ( .A(n97), .Q(n859) );
  NOR24 U473 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND23 U475 ( .A(B[20]), .B(A[20]), .Q(n145) );
  NAND22 U476 ( .A(n258), .B(n250), .Q(n248) );
  CLKIN3 U477 ( .A(n247), .Q(n886) );
  NAND24 U478 ( .A(n852), .B(n884), .Q(n422) );
  NOR23 U479 ( .A(n212), .B(n205), .Q(n203) );
  NOR24 U480 ( .A(n113), .B(n151), .Q(n111) );
  OAI212 U481 ( .A(n879), .B(n843), .C(n877), .Q(n164) );
  OAI212 U482 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  AOI212 U486 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR24 U488 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR24 U489 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND22 U490 ( .A(B[19]), .B(A[19]), .Q(n156) );
  XNR22 U491 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NAND24 U492 ( .A(n422), .B(n65), .Q(n63) );
  XNR22 U493 ( .A(n8), .B(n52), .Q(SUM[30]) );
  OAI211 U495 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  NAND21 U496 ( .A(A[8]), .B(B[8]), .Q(n245) );
  OAI211 U497 ( .A(n46), .B(n516), .C(n47), .Q(n45) );
  NAND24 U498 ( .A(n59), .B(n845), .Q(n46) );
  NOR23 U499 ( .A(n61), .B(n70), .Q(n59) );
  OAI212 U500 ( .A(n107), .B(n99), .C(n100), .Q(n674) );
  NOR23 U501 ( .A(B[20]), .B(A[20]), .Q(n144) );
  OAI212 U504 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI211 U505 ( .A(n213), .B(n205), .C(n206), .Q(n425) );
  INV1 U506 ( .A(n213), .Q(n900) );
  OAI212 U507 ( .A(n843), .B(n42), .C(n43), .Q(n41) );
  BUF15 U508 ( .A(n178), .Q(n843) );
  NOR24 U509 ( .A(B[23]), .B(A[23]), .Q(n117) );
  OAI210 U510 ( .A(n177), .B(n173), .C(n174), .Q(n756) );
  NAND22 U511 ( .A(A[21]), .B(B[21]), .Q(n138) );
  OAI212 U512 ( .A(n843), .B(n82), .C(n83), .Q(n81) );
  XNR22 U513 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NOR23 U514 ( .A(n70), .B(n6), .Q(n66) );
  NOR23 U515 ( .A(B[28]), .B(A[28]), .Q(n70) );
  INV1 U516 ( .A(n144), .Q(n881) );
  NAND21 U517 ( .A(A[23]), .B(B[23]), .Q(n118) );
  INV0 U519 ( .A(n155), .Q(n882) );
  NOR24 U520 ( .A(A[21]), .B(B[21]), .Q(n137) );
  NOR24 U521 ( .A(A[27]), .B(B[27]), .Q(n79) );
  OAI211 U522 ( .A(n126), .B(n870), .C(n127), .Q(n123) );
  INV1 U523 ( .A(n137), .Q(n871) );
  NOR24 U524 ( .A(n137), .B(n144), .Q(n135) );
  NOR24 U525 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND26 U526 ( .A(n97), .B(n423), .Q(n6) );
  NAND22 U527 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND22 U528 ( .A(A[18]), .B(B[18]), .Q(n163) );
  OAI212 U529 ( .A(n79), .B(n89), .C(n80), .Q(n78) );
  NOR24 U530 ( .A(n79), .B(n88), .Q(n423) );
  INV2 U531 ( .A(n88), .Q(n857) );
  NOR24 U532 ( .A(n106), .B(n99), .Q(n97) );
  NAND22 U533 ( .A(A[27]), .B(B[27]), .Q(n80) );
  INV2 U534 ( .A(n145), .Q(n880) );
  NAND20 U535 ( .A(n876), .B(n135), .Q(n129) );
  NAND23 U536 ( .A(n507), .B(n71), .Q(n67) );
  NAND22 U537 ( .A(n851), .B(n71), .Q(n10) );
  NAND21 U538 ( .A(n881), .B(n145), .Q(n18) );
  NAND21 U539 ( .A(n111), .B(n97), .Q(n91) );
  INV3 U540 ( .A(n135), .Q(n872) );
  AOI212 U541 ( .A(n98), .B(n423), .C(n78), .Q(n5) );
  AOI212 U543 ( .A(n674), .B(n423), .C(n78), .Q(n516) );
  NOR22 U544 ( .A(B[16]), .B(A[16]), .Q(n176) );
  INV3 U545 ( .A(n59), .Q(n850) );
  NAND21 U546 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND21 U547 ( .A(n876), .B(n122), .Q(n120) );
  NAND21 U548 ( .A(A[7]), .B(B[7]), .Q(n253) );
  CLKIN0 U549 ( .A(n173), .Q(n878) );
  NAND21 U550 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NOR22 U551 ( .A(B[7]), .B(A[7]), .Q(n252) );
  AOI210 U552 ( .A(n906), .B(n258), .C(n259), .Q(n257) );
  INV2 U553 ( .A(n51), .Q(n846) );
  INV0 U554 ( .A(n212), .Q(n901) );
  NAND21 U555 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND20 U556 ( .A(n896), .B(n253), .Q(n31) );
  INV2 U557 ( .A(n64), .Q(n852) );
  AOI212 U558 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  INV0 U559 ( .A(n171), .Q(n879) );
  INV0 U560 ( .A(n239), .Q(n894) );
  INV0 U561 ( .A(n107), .Q(n860) );
  AOI211 U562 ( .A(n756), .B(n875), .C(n873), .Q(n159) );
  INV0 U563 ( .A(n230), .Q(n890) );
  INV0 U564 ( .A(n244), .Q(n893) );
  INV0 U565 ( .A(n255), .Q(n887) );
  NOR22 U566 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NAND21 U567 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND20 U568 ( .A(A[9]), .B(B[9]), .Q(n242) );
  INV2 U569 ( .A(n39), .Q(n844) );
  INV3 U570 ( .A(n53), .Q(n849) );
  INV3 U571 ( .A(n219), .Q(n891) );
  INV3 U572 ( .A(n756), .Q(n877) );
  INV0 U573 ( .A(n240), .Q(n892) );
  INV3 U574 ( .A(n268), .Q(n906) );
  AOI211 U575 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U576 ( .A(n252), .B(n255), .Q(n250) );
  NOR21 U577 ( .A(n241), .B(n244), .Q(n239) );
  NOR21 U578 ( .A(n88), .B(n859), .Q(n84) );
  NOR21 U579 ( .A(n592), .B(n880), .Q(n141) );
  NAND20 U580 ( .A(n171), .B(n875), .Q(n158) );
  NAND22 U581 ( .A(n891), .B(n901), .Q(n208) );
  AOI211 U582 ( .A(n889), .B(n901), .C(n900), .Q(n209) );
  NAND22 U583 ( .A(n891), .B(n190), .Q(n188) );
  AOI211 U584 ( .A(n889), .B(n190), .C(n191), .Q(n189) );
  NAND20 U585 ( .A(n239), .B(n890), .Q(n226) );
  AOI210 U586 ( .A(n240), .B(n890), .C(n888), .Q(n227) );
  INV3 U587 ( .A(n231), .Q(n888) );
  INV3 U588 ( .A(n425), .Q(n897) );
  NOR20 U589 ( .A(n152), .B(n144), .Q(n592) );
  NAND22 U590 ( .A(n854), .B(n80), .Q(n11) );
  INV3 U591 ( .A(n79), .Q(n854) );
  NAND22 U592 ( .A(n853), .B(n851), .Q(n507) );
  INV3 U593 ( .A(n127), .Q(n868) );
  INV3 U594 ( .A(n126), .Q(n869) );
  INV3 U595 ( .A(n99), .Q(n862) );
  INV3 U596 ( .A(n61), .Q(n848) );
  INV3 U597 ( .A(n176), .Q(n883) );
  INV3 U598 ( .A(n274), .Q(n905) );
  NAND22 U599 ( .A(n904), .B(n261), .Q(n33) );
  INV3 U600 ( .A(n260), .Q(n904) );
  INV3 U601 ( .A(n265), .Q(n907) );
  INV3 U602 ( .A(n241), .Q(n895) );
  INV3 U603 ( .A(n252), .Q(n896) );
  NAND22 U604 ( .A(n909), .B(n272), .Q(n35) );
  INV3 U605 ( .A(n271), .Q(n909) );
  AOI211 U606 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U607 ( .A(n271), .B(n274), .Q(n269) );
  NOR21 U608 ( .A(n260), .B(n265), .Q(n258) );
  INV3 U609 ( .A(n277), .Q(n911) );
  INV3 U610 ( .A(n278), .Q(n913) );
  INV3 U611 ( .A(n266), .Q(n908) );
  NOR21 U612 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U613 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U614 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR21 U615 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR21 U616 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND22 U617 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND22 U618 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV3 U619 ( .A(n50), .Q(n845) );
  NOR21 U620 ( .A(A[30]), .B(B[30]), .Q(n50) );
  NOR21 U621 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR21 U622 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U623 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U624 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U625 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U626 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U627 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U628 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND22 U629 ( .A(A[0]), .B(B[0]), .Q(n281) );
  INV3 U630 ( .A(n280), .Q(n912) );
  NOR21 U631 ( .A(B[0]), .B(A[0]), .Q(n280) );
  XOR21 U632 ( .A(n30), .B(n886), .Q(SUM[8]) );
  NAND20 U633 ( .A(n893), .B(n245), .Q(n30) );
  XOR21 U634 ( .A(n36), .B(n911), .Q(SUM[2]) );
  NAND22 U635 ( .A(n905), .B(n275), .Q(n36) );
  XNR21 U636 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U637 ( .A(n895), .B(n242), .Q(n29) );
  XNR21 U638 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XOR20 U639 ( .A(n22), .B(n843), .Q(SUM[16]) );
  NAND20 U640 ( .A(n883), .B(n177), .Q(n22) );
  NAND20 U641 ( .A(n857), .B(n89), .Q(n12) );
  NAND20 U642 ( .A(n862), .B(n100), .Q(n13) );
  NAND22 U643 ( .A(n844), .B(n40), .Q(n7) );
  XNR21 U644 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NAND22 U645 ( .A(n174), .B(n878), .Q(n21) );
  NAND20 U646 ( .A(n858), .B(n107), .Q(n14) );
  XNR21 U647 ( .A(n18), .B(n146), .Q(SUM[20]) );
  XNR21 U648 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND20 U649 ( .A(n869), .B(n127), .Q(n16) );
  NAND20 U650 ( .A(n871), .B(n138), .Q(n17) );
  XNR21 U651 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND20 U652 ( .A(n865), .B(n118), .Q(n15) );
  NAND20 U653 ( .A(n163), .B(n875), .Q(n20) );
  NAND20 U654 ( .A(n156), .B(n882), .Q(n19) );
  XNR21 U655 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U656 ( .A(n901), .B(n213), .Q(n26) );
  XNR21 U657 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U658 ( .A(n206), .B(n898), .Q(n25) );
  XNR21 U659 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U660 ( .A(n902), .B(n195), .Q(n24) );
  XNR21 U661 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U662 ( .A(n885), .B(n186), .Q(n23) );
  NAND20 U663 ( .A(n848), .B(n62), .Q(n9) );
  XNR21 U664 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U666 ( .A(n890), .B(n231), .Q(n28) );
  XNR21 U667 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U668 ( .A(n903), .B(n224), .Q(n27) );
  XOR21 U669 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND22 U670 ( .A(n887), .B(n256), .Q(n32) );
  XOR21 U671 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U672 ( .A(n906), .B(n907), .C(n908), .Q(n262) );
  XNR21 U673 ( .A(n34), .B(n906), .Q(SUM[4]) );
  NAND22 U674 ( .A(n907), .B(n266), .Q(n34) );
  XNR21 U675 ( .A(n35), .B(n273), .Q(SUM[3]) );
  INV3 U676 ( .A(n38), .Q(SUM[0]) );
  NAND22 U677 ( .A(n912), .B(n281), .Q(n38) );
  XOR21 U678 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U679 ( .A(n913), .B(n279), .Q(n37) );
  INV3 U680 ( .A(n98), .Q(n861) );
endmodule


module adder_34 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_34_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_33_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n50,
         n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n416, n419, n486,
         n491, n492, n559, n563, n564, n637, n638, n643, n644, n717, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n869,
         n870, n871;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n802), .C(n121), .Q(n119) );
  OAI212 U127 ( .A(n129), .B(n801), .C(n130), .Q(n128) );
  OAI212 U141 ( .A(n140), .B(n802), .C(n141), .Q(n139) );
  OAI212 U165 ( .A(n158), .B(n801), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n844), .B(n801), .C(n845), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U197 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U233 ( .A(n208), .B(n826), .C(n209), .Q(n207) );
  OAI212 U257 ( .A(n226), .B(n826), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n840), .B(n826), .C(n838), .Q(n232) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n870), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U399 ( .A(n91), .B(n802), .C(n92), .Q(n90) );
  OAI212 U410 ( .A(n820), .B(n801), .C(n821), .Q(n108) );
  OAI212 U351 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U374 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  AOI212 U359 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  AOI212 U391 ( .A(n172), .B(n153), .C(n154), .Q(n486) );
  OAI212 U460 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U469 ( .A(n197), .B(n826), .C(n198), .Q(n196) );
  OAI212 U396 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U448 ( .A(n151), .B(n802), .C(n486), .Q(n146) );
  AOI212 U379 ( .A(n637), .B(n221), .C(n638), .Q(n559) );
  OAI212 U380 ( .A(n82), .B(n801), .C(n83), .Q(n81) );
  OAI212 U479 ( .A(n241), .B(n245), .C(n242), .Q(n416) );
  OAI212 U481 ( .A(n113), .B(n486), .C(n114), .Q(n419) );
  OAI212 U390 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U395 ( .A(n188), .B(n826), .C(n189), .Q(n187) );
  OAI212 U437 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI212 U456 ( .A(n126), .B(n831), .C(n127), .Q(n123) );
  OAI212 U377 ( .A(n64), .B(n802), .C(n65), .Q(n63) );
  OAI212 U387 ( .A(n73), .B(n802), .C(n74), .Q(n72) );
  OAI212 U398 ( .A(n102), .B(n801), .C(n103), .Q(n101) );
  OAI212 U430 ( .A(n799), .B(n155), .C(n156), .Q(n154) );
  OAI212 U453 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U465 ( .A(n223), .B(n231), .C(n224), .Q(n222) );
  AOI212 U468 ( .A(n416), .B(n221), .C(n222), .Q(n220) );
  OAI212 U394 ( .A(n244), .B(n826), .C(n245), .Q(n243) );
  OAI212 U475 ( .A(n53), .B(n802), .C(n54), .Q(n52) );
  OAI212 U476 ( .A(n42), .B(n802), .C(n43), .Q(n41) );
  OAI212 U509 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  XOR22 U349 ( .A(n717), .B(n214), .Q(SUM[12]) );
  INV3 U350 ( .A(n135), .Q(n833) );
  NAND22 U352 ( .A(A[20]), .B(B[20]), .Q(n145) );
  OAI210 U353 ( .A(n194), .B(n856), .C(n195), .Q(n191) );
  INV2 U354 ( .A(n204), .Q(n856) );
  OAI212 U355 ( .A(n223), .B(n231), .C(n224), .Q(n638) );
  NAND23 U356 ( .A(n563), .B(n564), .Q(SUM[17]) );
  NOR23 U357 ( .A(A[15]), .B(B[15]), .Q(n185) );
  CLKIN6 U358 ( .A(n857), .Q(n796) );
  AOI211 U360 ( .A(n112), .B(n55), .C(n56), .Q(n54) );
  NOR22 U361 ( .A(n807), .B(n6), .Q(n55) );
  OAI211 U362 ( .A(n807), .B(n5), .C(n808), .Q(n56) );
  XNR22 U363 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND21 U364 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NOR24 U365 ( .A(A[14]), .B(B[14]), .Q(n194) );
  BUF6 U366 ( .A(n88), .Q(n791) );
  XNR22 U367 ( .A(n16), .B(n128), .Q(SUM[22]) );
  INV3 U368 ( .A(n97), .Q(n815) );
  NAND22 U369 ( .A(n97), .B(n77), .Q(n6) );
  INV3 U370 ( .A(n151), .Q(n835) );
  INV0 U371 ( .A(n213), .Q(n862) );
  NOR21 U372 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND24 U373 ( .A(n171), .B(n153), .Q(n151) );
  NOR22 U375 ( .A(B[22]), .B(A[22]), .Q(n126) );
  INV3 U376 ( .A(n175), .Q(n825) );
  XNR21 U378 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U381 ( .A(n824), .B(n854), .Q(n644) );
  NOR22 U382 ( .A(n185), .B(n194), .Q(n183) );
  NOR22 U383 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR22 U384 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR21 U385 ( .A(n173), .B(n176), .Q(n171) );
  AOI211 U386 ( .A(n112), .B(n818), .C(n817), .Q(n103) );
  AOI211 U388 ( .A(n419), .B(n84), .C(n85), .Q(n83) );
  INV3 U389 ( .A(n139), .Q(n824) );
  NAND22 U392 ( .A(B[10]), .B(A[10]), .Q(n231) );
  XNR21 U393 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XNR21 U397 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND22 U400 ( .A(n491), .B(n492), .Q(SUM[16]) );
  NOR24 U401 ( .A(n212), .B(n796), .Q(n203) );
  NAND22 U402 ( .A(n797), .B(n21), .Q(n563) );
  NOR22 U403 ( .A(n117), .B(n126), .Q(n115) );
  NAND22 U404 ( .A(n19), .B(n157), .Q(n794) );
  NAND24 U405 ( .A(n792), .B(n793), .Q(n795) );
  NAND26 U406 ( .A(n794), .B(n795), .Q(SUM[19]) );
  INV3 U407 ( .A(n19), .Q(n792) );
  CLKIN6 U408 ( .A(n157), .Q(n793) );
  NAND20 U409 ( .A(n834), .B(n156), .Q(n19) );
  NOR23 U411 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NAND21 U412 ( .A(A[18]), .B(B[18]), .Q(n163) );
  CLKIN3 U413 ( .A(n230), .Q(n849) );
  NOR24 U414 ( .A(n223), .B(n230), .Q(n221) );
  NOR21 U415 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND21 U416 ( .A(n814), .B(n100), .Q(n13) );
  OAI212 U417 ( .A(n241), .B(n245), .C(n242), .Q(n637) );
  OAI211 U418 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  INV0 U419 ( .A(n241), .Q(n839) );
  CLKIN3 U420 ( .A(n231), .Q(n848) );
  NOR22 U421 ( .A(A[10]), .B(B[10]), .Q(n230) );
  AOI211 U422 ( .A(n112), .B(n66), .C(n67), .Q(n65) );
  INV6 U423 ( .A(n559), .Q(n837) );
  OAI211 U424 ( .A(n219), .B(n826), .C(n559), .Q(n214) );
  NAND22 U425 ( .A(n59), .B(n805), .Q(n46) );
  NOR22 U426 ( .A(n181), .B(n219), .Q(n179) );
  NAND23 U427 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR20 U428 ( .A(B[3]), .B(A[3]), .Q(n271) );
  CLKIN0 U429 ( .A(n212), .Q(n861) );
  NAND23 U431 ( .A(n203), .B(n183), .Q(n181) );
  NAND24 U432 ( .A(n643), .B(n644), .Q(SUM[21]) );
  NAND21 U433 ( .A(n111), .B(n55), .Q(n53) );
  NOR22 U434 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND20 U435 ( .A(n224), .B(n859), .Q(n27) );
  CLKIN6 U436 ( .A(n205), .Q(n857) );
  INV10 U438 ( .A(n800), .Q(n801) );
  XNR22 U439 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NAND21 U440 ( .A(B[13]), .B(A[13]), .Q(n206) );
  NOR23 U441 ( .A(A[13]), .B(B[13]), .Q(n205) );
  AOI212 U442 ( .A(n183), .B(n204), .C(n184), .Q(n182) );
  OAI211 U443 ( .A(n176), .B(n802), .C(n177), .Q(n797) );
  NAND21 U444 ( .A(A[26]), .B(B[26]), .Q(n89) );
  XNR22 U445 ( .A(n10), .B(n72), .Q(SUM[28]) );
  INV15 U446 ( .A(n800), .Q(n802) );
  NOR23 U447 ( .A(n194), .B(n858), .Q(n190) );
  NAND22 U449 ( .A(B[14]), .B(A[14]), .Q(n195) );
  OAI212 U450 ( .A(n185), .B(n195), .C(n186), .Q(n184) );
  NOR22 U451 ( .A(n79), .B(n791), .Q(n77) );
  NOR22 U452 ( .A(B[20]), .B(A[20]), .Q(n144) );
  AOI211 U454 ( .A(n836), .B(n122), .C(n123), .Q(n121) );
  XNR22 U455 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U457 ( .A(n813), .B(n89), .Q(n12) );
  OAI211 U458 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NAND22 U459 ( .A(B[9]), .B(A[9]), .Q(n242) );
  NAND21 U461 ( .A(A[21]), .B(B[21]), .Q(n138) );
  XNR22 U462 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NOR24 U463 ( .A(B[11]), .B(A[11]), .Q(n223) );
  XNR22 U464 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NOR23 U466 ( .A(n155), .B(n162), .Q(n153) );
  NOR22 U467 ( .A(B[12]), .B(A[12]), .Q(n212) );
  XNR22 U470 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NOR22 U471 ( .A(n99), .B(n106), .Q(n97) );
  INV0 U472 ( .A(n99), .Q(n814) );
  NAND22 U473 ( .A(n111), .B(n97), .Q(n91) );
  AOI211 U474 ( .A(n112), .B(n97), .C(n98), .Q(n92) );
  INV0 U477 ( .A(n194), .Q(n822) );
  NAND22 U478 ( .A(n865), .B(n802), .Q(n492) );
  NAND21 U480 ( .A(n867), .B(n186), .Q(n23) );
  INV0 U482 ( .A(n858), .Q(n798) );
  NAND22 U483 ( .A(A[12]), .B(B[12]), .Q(n213) );
  CLKIN1 U484 ( .A(n203), .Q(n858) );
  NAND20 U485 ( .A(n841), .B(n798), .Q(n197) );
  NOR21 U486 ( .A(B[24]), .B(A[24]), .Q(n106) );
  XNR22 U487 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NAND21 U488 ( .A(B[11]), .B(A[11]), .Q(n224) );
  OAI210 U489 ( .A(n791), .B(n816), .C(n89), .Q(n85) );
  OAI212 U490 ( .A(n176), .B(n802), .C(n177), .Q(n175) );
  XNR22 U491 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND22 U492 ( .A(A[16]), .B(B[16]), .Q(n177) );
  AOI211 U493 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  NAND21 U494 ( .A(A[24]), .B(B[24]), .Q(n107) );
  XNR22 U495 ( .A(n11), .B(n81), .Q(SUM[27]) );
  INV2 U496 ( .A(n106), .Q(n818) );
  NAND22 U497 ( .A(n835), .B(n122), .Q(n120) );
  INV6 U498 ( .A(n178), .Q(n800) );
  OAI212 U499 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  BUF6 U500 ( .A(n163), .Q(n799) );
  NAND22 U501 ( .A(n111), .B(n818), .Q(n102) );
  CLKIN3 U502 ( .A(n111), .Q(n820) );
  NAND22 U503 ( .A(n111), .B(n84), .Q(n82) );
  NAND22 U504 ( .A(n111), .B(n66), .Q(n64) );
  NOR24 U505 ( .A(n113), .B(n151), .Q(n111) );
  XNR22 U506 ( .A(n12), .B(n90), .Q(SUM[26]) );
  INV1 U507 ( .A(n6), .Q(n811) );
  AOI211 U508 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NOR22 U510 ( .A(B[23]), .B(A[23]), .Q(n117) );
  CLKIN1 U511 ( .A(n240), .Q(n838) );
  NAND20 U512 ( .A(A[19]), .B(B[19]), .Q(n156) );
  INV2 U513 ( .A(n802), .Q(n823) );
  NAND21 U514 ( .A(n809), .B(n71), .Q(n10) );
  NAND20 U515 ( .A(n851), .B(n799), .Q(n20) );
  OAI210 U516 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND20 U517 ( .A(n849), .B(n231), .Q(n28) );
  NAND21 U518 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NOR21 U519 ( .A(B[27]), .B(A[27]), .Q(n79) );
  AOI211 U520 ( .A(n419), .B(n811), .C(n812), .Q(n74) );
  INV1 U521 ( .A(n5), .Q(n812) );
  CLKIN0 U522 ( .A(n137), .Q(n855) );
  NOR21 U523 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR20 U524 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U525 ( .A(n486), .Q(n836) );
  AOI210 U526 ( .A(n837), .B(n203), .C(n204), .Q(n198) );
  NOR20 U527 ( .A(n46), .B(n6), .Q(n44) );
  NAND20 U528 ( .A(n171), .B(n851), .Q(n158) );
  CLKIN3 U529 ( .A(n59), .Q(n807) );
  NAND20 U530 ( .A(n239), .B(n221), .Q(n219) );
  NAND20 U531 ( .A(n841), .B(n190), .Q(n188) );
  NAND20 U532 ( .A(n841), .B(n861), .Q(n208) );
  NAND20 U533 ( .A(n239), .B(n849), .Q(n226) );
  NOR22 U534 ( .A(n137), .B(n144), .Q(n135) );
  NAND20 U535 ( .A(n832), .B(n145), .Q(n18) );
  NAND20 U536 ( .A(n818), .B(n107), .Q(n14) );
  CLKIN0 U537 ( .A(n171), .Q(n844) );
  INV0 U538 ( .A(n61), .Q(n806) );
  INV0 U539 ( .A(n70), .Q(n809) );
  NOR20 U540 ( .A(n212), .B(n862), .Q(n717) );
  NOR20 U541 ( .A(n241), .B(n244), .Q(n239) );
  NOR20 U542 ( .A(n252), .B(n255), .Q(n250) );
  NAND20 U543 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND20 U544 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U545 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U546 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U547 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U548 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NOR20 U549 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND20 U550 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U551 ( .A(n111), .B(n811), .Q(n73) );
  NAND20 U552 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U553 ( .A(n219), .Q(n841) );
  AOI211 U554 ( .A(n836), .B(n135), .C(n136), .Q(n130) );
  NAND22 U555 ( .A(n842), .B(n825), .Q(n564) );
  INV3 U556 ( .A(n21), .Q(n842) );
  AOI211 U557 ( .A(n837), .B(n861), .C(n862), .Q(n209) );
  INV3 U558 ( .A(n60), .Q(n808) );
  NAND22 U559 ( .A(n135), .B(n115), .Q(n113) );
  NAND22 U560 ( .A(n139), .B(n17), .Q(n643) );
  INV3 U561 ( .A(n17), .Q(n854) );
  NAND22 U562 ( .A(n22), .B(n823), .Q(n491) );
  INV3 U563 ( .A(n22), .Q(n865) );
  NAND22 U564 ( .A(n835), .B(n135), .Q(n129) );
  INV0 U565 ( .A(n172), .Q(n845) );
  AOI211 U566 ( .A(n846), .B(n258), .C(n259), .Q(n257) );
  INV3 U567 ( .A(n247), .Q(n826) );
  INV3 U568 ( .A(n268), .Q(n846) );
  INV3 U569 ( .A(n277), .Q(n870) );
  NAND22 U570 ( .A(n835), .B(n832), .Q(n140) );
  AOI211 U571 ( .A(n836), .B(n832), .C(n830), .Q(n141) );
  INV3 U572 ( .A(n145), .Q(n830) );
  NAND20 U573 ( .A(n857), .B(n206), .Q(n25) );
  NAND22 U574 ( .A(n819), .B(n118), .Q(n15) );
  INV3 U575 ( .A(n117), .Q(n819) );
  XOR21 U576 ( .A(n36), .B(n870), .Q(SUM[2]) );
  NAND22 U577 ( .A(n847), .B(n275), .Q(n36) );
  INV3 U578 ( .A(n274), .Q(n847) );
  XOR21 U579 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND22 U580 ( .A(n828), .B(n256), .Q(n32) );
  INV3 U581 ( .A(n255), .Q(n828) );
  XOR21 U582 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U583 ( .A(n846), .B(n864), .C(n863), .Q(n262) );
  NAND22 U584 ( .A(n829), .B(n261), .Q(n33) );
  INV3 U585 ( .A(n266), .Q(n863) );
  AOI211 U586 ( .A(n60), .B(n805), .C(n804), .Q(n47) );
  INV3 U587 ( .A(n51), .Q(n804) );
  NAND22 U588 ( .A(n810), .B(n80), .Q(n11) );
  INV3 U589 ( .A(n79), .Q(n810) );
  NAND22 U590 ( .A(n805), .B(n51), .Q(n8) );
  NAND22 U591 ( .A(n852), .B(n127), .Q(n16) );
  INV3 U592 ( .A(n126), .Q(n852) );
  XNR21 U593 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND22 U594 ( .A(n806), .B(n62), .Q(n9) );
  INV3 U595 ( .A(n791), .Q(n813) );
  INV3 U596 ( .A(n155), .Q(n834) );
  XNR21 U597 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND22 U598 ( .A(n839), .B(n242), .Q(n29) );
  NAND22 U599 ( .A(n822), .B(n195), .Q(n24) );
  XNR21 U600 ( .A(n28), .B(n232), .Q(SUM[10]) );
  INV3 U601 ( .A(n239), .Q(n840) );
  XNR21 U602 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND22 U603 ( .A(n827), .B(n253), .Q(n31) );
  INV3 U604 ( .A(n252), .Q(n827) );
  NOR21 U605 ( .A(n61), .B(n70), .Q(n59) );
  NOR21 U606 ( .A(n126), .B(n833), .Q(n122) );
  NOR21 U607 ( .A(n791), .B(n815), .Q(n84) );
  NOR21 U608 ( .A(n70), .B(n6), .Q(n66) );
  NAND22 U609 ( .A(n855), .B(n138), .Q(n17) );
  INV0 U610 ( .A(n185), .Q(n867) );
  AOI210 U611 ( .A(n172), .B(n851), .C(n850), .Q(n159) );
  INV3 U612 ( .A(n799), .Q(n850) );
  NAND21 U613 ( .A(n174), .B(n843), .Q(n21) );
  INV0 U614 ( .A(n173), .Q(n843) );
  NAND22 U615 ( .A(n866), .B(n177), .Q(n22) );
  INV3 U616 ( .A(n260), .Q(n829) );
  INV0 U617 ( .A(n98), .Q(n816) );
  INV2 U618 ( .A(n136), .Q(n831) );
  AOI211 U619 ( .A(n837), .B(n190), .C(n191), .Q(n189) );
  AOI211 U620 ( .A(n240), .B(n849), .C(n848), .Q(n227) );
  INV3 U621 ( .A(n107), .Q(n817) );
  INV3 U622 ( .A(n144), .Q(n832) );
  INV3 U623 ( .A(n162), .Q(n851) );
  XOR21 U624 ( .A(n30), .B(n826), .Q(SUM[8]) );
  NAND22 U625 ( .A(n860), .B(n245), .Q(n30) );
  INV2 U626 ( .A(n244), .Q(n860) );
  XNR21 U627 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U628 ( .A(n853), .B(n272), .Q(n35) );
  INV3 U629 ( .A(n271), .Q(n853) );
  INV3 U630 ( .A(n265), .Q(n864) );
  XNR21 U631 ( .A(n34), .B(n846), .Q(SUM[4]) );
  NAND22 U632 ( .A(n864), .B(n266), .Q(n34) );
  AOI211 U633 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U634 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U635 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U636 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  XOR21 U637 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U638 ( .A(n871), .B(n279), .Q(n37) );
  INV3 U639 ( .A(n278), .Q(n871) );
  NOR21 U640 ( .A(n260), .B(n265), .Q(n258) );
  NOR21 U641 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NAND22 U642 ( .A(n803), .B(n40), .Q(n7) );
  NAND22 U643 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR21 U644 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR20 U645 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV3 U646 ( .A(n50), .Q(n805) );
  INV3 U647 ( .A(n39), .Q(n803) );
  NAND20 U648 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND20 U649 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND20 U650 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND20 U651 ( .A(A[3]), .B(B[3]), .Q(n272) );
  INV3 U652 ( .A(n38), .Q(SUM[0]) );
  NAND22 U653 ( .A(n869), .B(n281), .Q(n38) );
  INV3 U654 ( .A(n280), .Q(n869) );
  NOR20 U655 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U656 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NOR20 U657 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND20 U658 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U659 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NOR20 U660 ( .A(B[2]), .B(A[2]), .Q(n274) );
  INV2 U661 ( .A(n223), .Q(n859) );
  NAND21 U662 ( .A(B[17]), .B(A[17]), .Q(n174) );
  NOR22 U663 ( .A(B[17]), .B(A[17]), .Q(n173) );
  INV3 U664 ( .A(n176), .Q(n866) );
  NOR22 U665 ( .A(B[16]), .B(A[16]), .Q(n176) );
  INV2 U666 ( .A(n419), .Q(n821) );
  AOI210 U667 ( .A(n419), .B(n44), .C(n45), .Q(n43) );
  NOR21 U668 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U669 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR21 U670 ( .A(B[5]), .B(A[5]), .Q(n260) );
endmodule


module adder_33 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_33_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n61, n62,
         n67, n68, n69, n70, n71, n74, n75, n76, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n95, n96, n97, n98, n99, n100, n105,
         n106, n107, n108, n109, n112, n113, n114, n115, n116, n121, n122,
         n123, n124, n125, n126, n127, n130, n131, n132, n136, n141, n142,
         n143, n144, n145, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n163, n164, n165, n166, n167, n168,
         n173, n174, n175, n176, n177, n180, n181, n182, n183, n184, n189,
         n190, n191, n192, n193, n194, n195, n198, n199, n200, n203, n204,
         n209, n210, n211, n212, n213, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n228, n229, n230, n231, n236, n237,
         n238, n241, n242, n244, n245, n246, n247, n248, n249, n250, n251,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n265, n266, n267, n268, n269, n405, n479, n481, n486, n551, n554,
         n555, n558, n559, n630, n631, n704, n705, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n849, n850, n851,
         n852, n853, n854, n855;

  OAI212 U74 ( .A(n88), .B(n785), .C(n89), .Q(n87) );
  OAI212 U94 ( .A(n113), .B(n105), .C(n106), .Q(n100) );
  OAI212 U100 ( .A(n108), .B(n785), .C(n109), .Q(n107) );
  OAI212 U134 ( .A(n481), .B(n785), .C(n828), .Q(n132) );
  OAI212 U142 ( .A(n145), .B(n141), .C(n142), .Q(n136) );
  AOI212 U154 ( .A(n405), .B(n147), .C(n148), .Q(n1) );
  OAI212 U186 ( .A(n181), .B(n173), .C(n174), .Q(n168) );
  OAI212 U247 ( .A(n216), .B(n244), .C(n217), .Q(n215) );
  OAI212 U290 ( .A(n251), .B(n247), .C(n248), .Q(n246) );
  OAI212 U296 ( .A(n250), .B(n851), .C(n251), .Q(n249) );
  OAI212 U303 ( .A(n254), .B(n256), .C(n255), .Q(n253) );
  OAI212 U311 ( .A(n263), .B(n259), .C(n260), .Q(n258) );
  OAI212 U317 ( .A(n262), .B(n850), .C(n263), .Q(n261) );
  OAI212 U324 ( .A(n269), .B(n266), .C(n267), .Q(n265) );
  OAI212 U403 ( .A(n97), .B(n785), .C(n98), .Q(n96) );
  OAI212 U356 ( .A(n216), .B(n244), .C(n217), .Q(n405) );
  OAI212 U388 ( .A(n176), .B(n821), .C(n177), .Q(n175) );
  OAI212 U415 ( .A(n799), .B(n785), .C(n797), .Q(n76) );
  OAI212 U419 ( .A(n184), .B(n149), .C(n150), .Q(n148) );
  OAI212 U427 ( .A(n199), .B(n191), .C(n192), .Q(n190) );
  OAI212 U380 ( .A(n57), .B(n47), .C(n48), .Q(n46) );
  OAI212 U433 ( .A(n194), .B(n821), .C(n195), .Q(n193) );
  AOI212 U343 ( .A(n136), .B(n121), .C(n122), .Q(n116) );
  OAI212 U410 ( .A(n70), .B(n785), .C(n71), .Q(n69) );
  OAI212 U401 ( .A(n39), .B(n785), .C(n40), .Q(n38) );
  OAI212 U352 ( .A(n115), .B(n785), .C(n116), .Q(n114) );
  OAI212 U374 ( .A(n212), .B(n821), .C(n213), .Q(n211) );
  OAI212 U466 ( .A(n75), .B(n67), .C(n68), .Q(n62) );
  OAI212 U469 ( .A(n54), .B(n793), .C(n57), .Q(n53) );
  OAI212 U484 ( .A(n156), .B(n821), .C(n157), .Q(n155) );
  OAI212 U337 ( .A(n126), .B(n785), .C(n127), .Q(n704) );
  OAI212 U348 ( .A(n59), .B(n785), .C(n60), .Q(n58) );
  OAI212 U338 ( .A(n126), .B(n785), .C(n127), .Q(n125) );
  OAI212 U461 ( .A(n225), .B(n835), .C(n228), .Q(n224) );
  AOI212 U339 ( .A(n2), .B(n52), .C(n53), .Q(n51) );
  NOR23 U340 ( .A(B[12]), .B(A[12]), .Q(n209) );
  XNR22 U341 ( .A(n21), .B(n193), .Q(SUM[14]) );
  XNR22 U342 ( .A(n11), .B(n107), .Q(SUM[24]) );
  XOR22 U344 ( .A(n24), .B(n821), .Q(SUM[11]) );
  CLKIN12 U345 ( .A(n215), .Q(n821) );
  NOR23 U346 ( .A(B[22]), .B(A[22]), .Q(n123) );
  OAI212 U347 ( .A(n236), .B(n242), .C(n237), .Q(n231) );
  NAND23 U349 ( .A(B[8]), .B(A[8]), .Q(n237) );
  NAND23 U350 ( .A(A[7]), .B(B[7]), .Q(n242) );
  OAI211 U351 ( .A(n50), .B(n785), .C(n51), .Q(n49) );
  NAND22 U353 ( .A(n3), .B(n52), .Q(n50) );
  NAND24 U354 ( .A(n630), .B(n631), .Q(SUM[22]) );
  NAND28 U355 ( .A(n167), .B(n151), .Q(n149) );
  NOR24 U357 ( .A(n153), .B(n160), .Q(n151) );
  NAND24 U358 ( .A(n781), .B(n782), .Q(n783) );
  NAND24 U359 ( .A(n783), .B(n210), .Q(n204) );
  INV4 U360 ( .A(n213), .Q(n781) );
  INV6 U361 ( .A(n209), .Q(n782) );
  NAND23 U362 ( .A(A[11]), .B(B[11]), .Q(n213) );
  OAI210 U363 ( .A(n95), .B(n85), .C(n86), .Q(n84) );
  NOR22 U364 ( .A(n85), .B(n92), .Q(n83) );
  NOR24 U365 ( .A(n191), .B(n198), .Q(n189) );
  NOR22 U366 ( .A(B[13]), .B(A[13]), .Q(n198) );
  XNR22 U367 ( .A(n18), .B(n164), .Q(SUM[17]) );
  INV3 U368 ( .A(n481), .Q(n826) );
  INV0 U369 ( .A(n130), .Q(n808) );
  INV3 U370 ( .A(n486), .Q(n833) );
  NOR21 U371 ( .A(B[21]), .B(A[21]), .Q(n130) );
  NOR21 U372 ( .A(n123), .B(n130), .Q(n121) );
  NOR21 U373 ( .A(B[23]), .B(A[23]), .Q(n112) );
  NOR22 U375 ( .A(n220), .B(n225), .Q(n218) );
  INV3 U376 ( .A(n144), .Q(n827) );
  NOR21 U377 ( .A(B[26]), .B(A[26]), .Q(n85) );
  NOR22 U378 ( .A(B[19]), .B(A[19]), .Q(n144) );
  INV3 U379 ( .A(n132), .Q(n814) );
  NOR23 U381 ( .A(A[10]), .B(B[10]), .Q(n220) );
  NOR22 U382 ( .A(B[11]), .B(A[11]), .Q(n212) );
  NAND26 U383 ( .A(n554), .B(n555), .Q(SUM[23]) );
  NAND24 U384 ( .A(n804), .B(n809), .Q(n555) );
  XOR21 U385 ( .A(n27), .B(n238), .Q(SUM[8]) );
  XNR21 U386 ( .A(n19), .B(n175), .Q(SUM[16]) );
  NOR23 U387 ( .A(B[18]), .B(A[18]), .Q(n153) );
  NAND22 U389 ( .A(n826), .B(n121), .Q(n115) );
  CLKIN3 U390 ( .A(n131), .Q(n811) );
  NAND21 U391 ( .A(n846), .B(n210), .Q(n23) );
  NAND21 U392 ( .A(A[12]), .B(B[12]), .Q(n210) );
  CLKIN6 U393 ( .A(n114), .Q(n809) );
  NAND23 U394 ( .A(n203), .B(n189), .Q(n183) );
  OAI212 U395 ( .A(n228), .B(n220), .C(n221), .Q(n219) );
  NOR24 U396 ( .A(A[8]), .B(B[8]), .Q(n236) );
  NAND23 U397 ( .A(n479), .B(n82), .Q(n2) );
  AOI211 U398 ( .A(n100), .B(n83), .C(n84), .Q(n82) );
  NOR22 U399 ( .A(B[20]), .B(A[20]), .Q(n141) );
  NAND26 U400 ( .A(n558), .B(n559), .Q(SUM[21]) );
  NOR24 U402 ( .A(B[16]), .B(A[16]), .Q(n173) );
  NAND21 U404 ( .A(n832), .B(n167), .Q(n165) );
  INV2 U405 ( .A(n183), .Q(n832) );
  XNR22 U406 ( .A(n23), .B(n211), .Q(SUM[12]) );
  NAND22 U407 ( .A(A[15]), .B(B[15]), .Q(n181) );
  NAND21 U408 ( .A(A[16]), .B(B[16]), .Q(n174) );
  OAI212 U409 ( .A(n163), .B(n153), .C(n154), .Q(n152) );
  XNR22 U411 ( .A(n22), .B(n200), .Q(SUM[13]) );
  OAI211 U412 ( .A(n840), .B(n821), .C(n838), .Q(n200) );
  NAND22 U413 ( .A(n784), .B(n805), .Q(n108) );
  OAI211 U414 ( .A(n236), .B(n242), .C(n237), .Q(n705) );
  NAND21 U416 ( .A(A[20]), .B(B[20]), .Q(n142) );
  NAND21 U417 ( .A(n845), .B(n154), .Q(n17) );
  XNR22 U418 ( .A(n4), .B(n38), .Q(SUM[31]) );
  NAND22 U420 ( .A(n844), .B(n242), .Q(n28) );
  NAND22 U421 ( .A(A[19]), .B(B[19]), .Q(n145) );
  XNR22 U422 ( .A(n5), .B(n49), .Q(SUM[30]) );
  OAI212 U423 ( .A(n183), .B(n821), .C(n486), .Q(n182) );
  AOI212 U424 ( .A(n204), .B(n189), .C(n190), .Q(n486) );
  XNR22 U425 ( .A(n6), .B(n58), .Q(SUM[29]) );
  BUF15 U426 ( .A(n1), .Q(n785) );
  NAND21 U428 ( .A(n826), .B(n808), .Q(n126) );
  NAND24 U429 ( .A(n807), .B(n814), .Q(n559) );
  AOI212 U430 ( .A(n189), .B(n204), .C(n190), .Q(n184) );
  AOI212 U431 ( .A(n168), .B(n151), .C(n152), .Q(n150) );
  AOI211 U432 ( .A(n815), .B(n168), .C(n813), .Q(n551) );
  NOR23 U434 ( .A(B[14]), .B(A[14]), .Q(n191) );
  NOR24 U435 ( .A(B[9]), .B(A[9]), .Q(n225) );
  AOI211 U436 ( .A(n833), .B(n167), .C(n168), .Q(n166) );
  NAND21 U437 ( .A(A[14]), .B(B[14]), .Q(n192) );
  XNR22 U438 ( .A(n17), .B(n155), .Q(SUM[18]) );
  NOR22 U439 ( .A(B[15]), .B(A[15]), .Q(n180) );
  NAND22 U440 ( .A(B[13]), .B(A[13]), .Q(n199) );
  NOR23 U441 ( .A(B[17]), .B(A[17]), .Q(n160) );
  NOR23 U442 ( .A(n173), .B(n180), .Q(n167) );
  NAND21 U443 ( .A(n784), .B(n99), .Q(n97) );
  INV3 U444 ( .A(n99), .Q(n801) );
  AOI211 U445 ( .A(n810), .B(n99), .C(n100), .Q(n98) );
  NOR22 U446 ( .A(n105), .B(n112), .Q(n99) );
  OAI212 U447 ( .A(n131), .B(n123), .C(n124), .Q(n122) );
  NAND21 U448 ( .A(A[22]), .B(B[22]), .Q(n124) );
  NOR22 U449 ( .A(B[25]), .B(A[25]), .Q(n92) );
  XOR22 U450 ( .A(n16), .B(n785), .Q(SUM[19]) );
  OAI212 U451 ( .A(n144), .B(n785), .C(n145), .Q(n143) );
  OAI211 U452 ( .A(n165), .B(n821), .C(n166), .Q(n164) );
  XNR22 U453 ( .A(n8), .B(n76), .Q(SUM[27]) );
  XNR22 U454 ( .A(n15), .B(n143), .Q(SUM[20]) );
  XNR22 U455 ( .A(n10), .B(n96), .Q(SUM[25]) );
  XNR22 U456 ( .A(n9), .B(n87), .Q(SUM[26]) );
  NAND21 U457 ( .A(A[10]), .B(B[10]), .Q(n221) );
  NAND20 U458 ( .A(n829), .B(n95), .Q(n10) );
  OAI211 U459 ( .A(n92), .B(n802), .C(n95), .Q(n91) );
  INV0 U460 ( .A(n220), .Q(n823) );
  NAND20 U462 ( .A(n230), .B(n218), .Q(n216) );
  NAND21 U463 ( .A(n815), .B(n163), .Q(n18) );
  INV2 U464 ( .A(n163), .Q(n813) );
  NAND21 U465 ( .A(A[17]), .B(B[17]), .Q(n163) );
  NAND21 U467 ( .A(A[21]), .B(B[21]), .Q(n131) );
  NAND21 U468 ( .A(n805), .B(n113), .Q(n12) );
  NAND22 U470 ( .A(A[23]), .B(B[23]), .Q(n113) );
  NOR22 U471 ( .A(n81), .B(n115), .Q(n3) );
  INV2 U472 ( .A(n209), .Q(n846) );
  NOR22 U473 ( .A(n209), .B(n212), .Q(n203) );
  XNR22 U474 ( .A(n7), .B(n69), .Q(SUM[28]) );
  NOR20 U475 ( .A(n47), .B(n54), .Q(n45) );
  NOR22 U476 ( .A(B[24]), .B(A[24]), .Q(n105) );
  NAND21 U477 ( .A(A[27]), .B(B[27]), .Q(n75) );
  NAND21 U478 ( .A(A[29]), .B(B[29]), .Q(n57) );
  NAND22 U479 ( .A(n798), .B(n810), .Q(n479) );
  INV0 U480 ( .A(n92), .Q(n829) );
  INV3 U481 ( .A(n115), .Q(n784) );
  CLKIN3 U482 ( .A(n705), .Q(n835) );
  INV0 U483 ( .A(n81), .Q(n798) );
  NAND22 U485 ( .A(n794), .B(n75), .Q(n8) );
  AOI211 U486 ( .A(n833), .B(n817), .C(n816), .Q(n177) );
  NAND20 U487 ( .A(A[25]), .B(B[25]), .Q(n95) );
  NOR22 U488 ( .A(B[28]), .B(A[28]), .Q(n67) );
  NAND20 U489 ( .A(A[18]), .B(B[18]), .Q(n154) );
  INV0 U490 ( .A(n212), .Q(n839) );
  AOI211 U491 ( .A(n2), .B(n794), .C(n795), .Q(n71) );
  NAND20 U492 ( .A(n841), .B(n174), .Q(n19) );
  NAND20 U493 ( .A(n847), .B(n192), .Q(n21) );
  CLKIN2 U494 ( .A(n3), .Q(n799) );
  INV0 U495 ( .A(n112), .Q(n805) );
  CLKIN0 U496 ( .A(n203), .Q(n840) );
  NAND20 U497 ( .A(n831), .B(n199), .Q(n22) );
  INV0 U498 ( .A(n225), .Q(n842) );
  NAND20 U499 ( .A(n3), .B(n788), .Q(n39) );
  NOR23 U500 ( .A(n149), .B(n183), .Q(n147) );
  INV3 U501 ( .A(n116), .Q(n810) );
  CLKIN3 U502 ( .A(n2), .Q(n797) );
  NAND20 U503 ( .A(n203), .B(n831), .Q(n194) );
  NAND20 U504 ( .A(n61), .B(n45), .Q(n43) );
  NAND20 U505 ( .A(n827), .B(n145), .Q(n16) );
  AOI211 U506 ( .A(n833), .B(n158), .C(n812), .Q(n157) );
  INV2 U507 ( .A(n551), .Q(n812) );
  AOI212 U508 ( .A(n218), .B(n231), .C(n219), .Q(n217) );
  CLKIN0 U509 ( .A(n167), .Q(n818) );
  NAND20 U510 ( .A(n817), .B(n181), .Q(n20) );
  INV0 U511 ( .A(n173), .Q(n841) );
  INV0 U512 ( .A(n191), .Q(n847) );
  NAND20 U513 ( .A(n142), .B(n830), .Q(n15) );
  NAND20 U514 ( .A(n791), .B(n68), .Q(n7) );
  INV0 U515 ( .A(n54), .Q(n790) );
  INV0 U516 ( .A(n85), .Q(n796) );
  CLKIN3 U517 ( .A(n61), .Q(n792) );
  NAND20 U518 ( .A(n842), .B(n228), .Q(n26) );
  INV0 U519 ( .A(n242), .Q(n843) );
  CLKIN1 U520 ( .A(n62), .Q(n793) );
  AOI210 U521 ( .A(n62), .B(n45), .C(n46), .Q(n44) );
  AOI210 U522 ( .A(n2), .B(n788), .C(n789), .Q(n40) );
  NAND20 U523 ( .A(n808), .B(n131), .Q(n14) );
  INV2 U524 ( .A(n241), .Q(n844) );
  INV1 U525 ( .A(n74), .Q(n794) );
  INV0 U526 ( .A(n236), .Q(n836) );
  NOR20 U527 ( .A(n236), .B(n241), .Q(n230) );
  NOR20 U528 ( .A(n247), .B(n250), .Q(n245) );
  NOR20 U529 ( .A(B[30]), .B(A[30]), .Q(n47) );
  NOR20 U530 ( .A(B[5]), .B(A[5]), .Q(n250) );
  NAND20 U531 ( .A(A[26]), .B(B[26]), .Q(n86) );
  NAND20 U532 ( .A(A[24]), .B(B[24]), .Q(n106) );
  NAND20 U533 ( .A(A[30]), .B(B[30]), .Q(n48) );
  INV0 U534 ( .A(n136), .Q(n828) );
  AOI211 U535 ( .A(n2), .B(n61), .C(n62), .Q(n60) );
  NAND22 U536 ( .A(n99), .B(n83), .Q(n81) );
  NAND22 U537 ( .A(n132), .B(n14), .Q(n558) );
  INV3 U538 ( .A(n14), .Q(n807) );
  NAND22 U539 ( .A(n13), .B(n125), .Q(n630) );
  NAND22 U540 ( .A(n824), .B(n806), .Q(n631) );
  NAND22 U541 ( .A(n830), .B(n827), .Q(n481) );
  NAND22 U542 ( .A(n114), .B(n12), .Q(n554) );
  INV3 U543 ( .A(n12), .Q(n804) );
  NAND22 U544 ( .A(n3), .B(n61), .Q(n59) );
  NAND21 U545 ( .A(n3), .B(n794), .Q(n70) );
  NAND22 U546 ( .A(n784), .B(n90), .Q(n88) );
  NAND22 U547 ( .A(n832), .B(n158), .Q(n156) );
  INV3 U548 ( .A(n704), .Q(n806) );
  NAND22 U549 ( .A(n832), .B(n817), .Q(n176) );
  INV0 U550 ( .A(n204), .Q(n838) );
  INV3 U551 ( .A(n13), .Q(n824) );
  INV3 U552 ( .A(n43), .Q(n788) );
  INV3 U553 ( .A(n244), .Q(n820) );
  INV3 U554 ( .A(n253), .Q(n851) );
  INV3 U555 ( .A(n265), .Q(n850) );
  AOI211 U556 ( .A(n820), .B(n844), .C(n843), .Q(n238) );
  NAND22 U557 ( .A(n836), .B(n237), .Q(n27) );
  XOR21 U558 ( .A(n25), .B(n222), .Q(SUM[10]) );
  NAND22 U559 ( .A(n823), .B(n221), .Q(n25) );
  AOI211 U560 ( .A(n820), .B(n223), .C(n224), .Q(n222) );
  NAND22 U561 ( .A(n796), .B(n86), .Q(n9) );
  INV3 U562 ( .A(n153), .Q(n845) );
  NAND22 U563 ( .A(n790), .B(n57), .Q(n6) );
  INV3 U564 ( .A(n67), .Q(n791) );
  XNR21 U565 ( .A(n28), .B(n820), .Q(SUM[7]) );
  XNR21 U566 ( .A(n29), .B(n249), .Q(SUM[6]) );
  NAND22 U567 ( .A(n819), .B(n248), .Q(n29) );
  INV3 U568 ( .A(n247), .Q(n819) );
  NAND22 U569 ( .A(n800), .B(n106), .Q(n11) );
  INV3 U570 ( .A(n105), .Q(n800) );
  NAND22 U571 ( .A(n787), .B(n48), .Q(n5) );
  INV3 U572 ( .A(n47), .Q(n787) );
  XOR21 U573 ( .A(n851), .B(n30), .Q(SUM[5]) );
  NAND22 U574 ( .A(n822), .B(n251), .Q(n30) );
  INV3 U575 ( .A(n250), .Q(n822) );
  NOR21 U576 ( .A(n67), .B(n74), .Q(n61) );
  NAND22 U577 ( .A(n839), .B(n213), .Q(n24) );
  INV3 U578 ( .A(n199), .Q(n834) );
  XNR21 U579 ( .A(n20), .B(n182), .Q(SUM[15]) );
  NOR21 U580 ( .A(n92), .B(n801), .Q(n90) );
  NOR21 U581 ( .A(n160), .B(n818), .Q(n158) );
  AOI210 U582 ( .A(n136), .B(n808), .C(n811), .Q(n127) );
  XOR21 U583 ( .A(n26), .B(n229), .Q(SUM[9]) );
  AOI211 U584 ( .A(n820), .B(n230), .C(n705), .Q(n229) );
  NAND22 U585 ( .A(n825), .B(n124), .Q(n13) );
  INV3 U586 ( .A(n123), .Q(n825) );
  AOI211 U587 ( .A(n810), .B(n90), .C(n91), .Q(n89) );
  INV3 U588 ( .A(n100), .Q(n802) );
  INV3 U589 ( .A(n75), .Q(n795) );
  AOI210 U590 ( .A(n810), .B(n805), .C(n803), .Q(n109) );
  INV3 U591 ( .A(n113), .Q(n803) );
  INV3 U592 ( .A(n181), .Q(n816) );
  INV3 U593 ( .A(n44), .Q(n789) );
  INV3 U594 ( .A(n180), .Q(n817) );
  INV3 U595 ( .A(n198), .Q(n831) );
  INV3 U596 ( .A(n141), .Q(n830) );
  INV3 U597 ( .A(n160), .Q(n815) );
  NOR21 U598 ( .A(n54), .B(n792), .Q(n52) );
  AOI211 U599 ( .A(n245), .B(n253), .C(n246), .Q(n244) );
  XOR21 U600 ( .A(n31), .B(n256), .Q(SUM[4]) );
  NAND22 U601 ( .A(n855), .B(n255), .Q(n31) );
  INV3 U602 ( .A(n254), .Q(n855) );
  XOR21 U603 ( .A(n33), .B(n850), .Q(SUM[2]) );
  NAND22 U604 ( .A(n853), .B(n263), .Q(n33) );
  INV3 U605 ( .A(n262), .Q(n853) );
  XOR21 U606 ( .A(n269), .B(n34), .Q(SUM[1]) );
  NAND22 U607 ( .A(n852), .B(n267), .Q(n34) );
  INV3 U608 ( .A(n266), .Q(n852) );
  XNR21 U609 ( .A(n32), .B(n261), .Q(SUM[3]) );
  NAND22 U610 ( .A(n854), .B(n260), .Q(n32) );
  INV3 U611 ( .A(n259), .Q(n854) );
  AOI211 U612 ( .A(n265), .B(n257), .C(n258), .Q(n256) );
  NOR21 U613 ( .A(n259), .B(n262), .Q(n257) );
  NOR21 U614 ( .A(n225), .B(n837), .Q(n223) );
  INV3 U615 ( .A(n230), .Q(n837) );
  NAND22 U616 ( .A(n786), .B(n37), .Q(n4) );
  NAND20 U617 ( .A(A[31]), .B(B[31]), .Q(n37) );
  NOR21 U618 ( .A(B[29]), .B(A[29]), .Q(n54) );
  NOR21 U619 ( .A(B[6]), .B(A[6]), .Q(n247) );
  NOR21 U620 ( .A(B[27]), .B(A[27]), .Q(n74) );
  NOR20 U621 ( .A(B[7]), .B(A[7]), .Q(n241) );
  NAND22 U622 ( .A(B[9]), .B(A[9]), .Q(n228) );
  NAND20 U623 ( .A(A[28]), .B(B[28]), .Q(n68) );
  INV3 U624 ( .A(n36), .Q(n786) );
  NOR20 U625 ( .A(B[31]), .B(A[31]), .Q(n36) );
  NAND20 U626 ( .A(A[5]), .B(B[5]), .Q(n251) );
  NAND20 U627 ( .A(A[6]), .B(B[6]), .Q(n248) );
  INV3 U628 ( .A(n35), .Q(SUM[0]) );
  NAND22 U629 ( .A(n849), .B(n269), .Q(n35) );
  INV3 U630 ( .A(n268), .Q(n849) );
  NOR20 U631 ( .A(B[0]), .B(A[0]), .Q(n268) );
  NOR20 U632 ( .A(B[3]), .B(A[3]), .Q(n259) );
  NOR20 U633 ( .A(B[2]), .B(A[2]), .Q(n262) );
  NAND20 U634 ( .A(A[0]), .B(B[0]), .Q(n269) );
  NAND20 U635 ( .A(A[2]), .B(B[2]), .Q(n263) );
  NOR20 U636 ( .A(B[1]), .B(A[1]), .Q(n266) );
  NOR20 U637 ( .A(B[4]), .B(A[4]), .Q(n254) );
  NAND20 U638 ( .A(A[1]), .B(B[1]), .Q(n267) );
  NAND20 U639 ( .A(A[3]), .B(B[3]), .Q(n260) );
  NAND20 U640 ( .A(A[4]), .B(B[4]), .Q(n255) );
  AOI210 U641 ( .A(n204), .B(n831), .C(n834), .Q(n195) );
endmodule


module adder_32 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_32_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module reg_9 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30,
         n32, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n109, n110, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395;

  DF3 Dout_reg_16_ ( .D(n88), .C(Clk), .Q(Dout[16]), .QN(n87) );
  DF3 Dout_reg_14_ ( .D(n90), .C(Clk), .Q(Dout[14]), .QN(n73) );
  DF3 Dout_reg_13_ ( .D(n91), .C(Clk), .Q(Dout[13]), .QN(n72) );
  DF3 Dout_reg_12_ ( .D(n92), .C(Clk), .Q(Dout[12]), .QN(n71) );
  DF3 Dout_reg_11_ ( .D(n93), .C(Clk), .Q(Dout[11]), .QN(n81) );
  DF3 Dout_reg_10_ ( .D(n94), .C(Clk), .Q(Dout[10]), .QN(n80) );
  DF3 Dout_reg_8_ ( .D(n96), .C(Clk), .Q(Dout[8]), .QN(n78) );
  DF3 Dout_reg_7_ ( .D(n97), .C(Clk), .Q(Dout[7]), .QN(n77) );
  DF3 Dout_reg_6_ ( .D(n98), .C(Clk), .Q(Dout[6]), .QN(n76) );
  DF3 Dout_reg_5_ ( .D(n99), .C(Clk), .Q(Dout[5]), .QN(n82) );
  DF3 Dout_reg_4_ ( .D(n100), .C(Clk), .Q(Dout[4]), .QN(n85) );
  DF3 Dout_reg_2_ ( .D(n102), .C(Clk), .Q(Dout[2]), .QN(n75) );
  DF3 Dout_reg_0_ ( .D(n104), .C(Clk), .Q(Dout[0]), .QN(n86) );
  DF3 Dout_reg_15_ ( .D(n89), .C(Clk), .Q(Dout[15]), .QN(n74) );
  DF3 Dout_reg_3_ ( .D(n101), .C(Clk), .Q(Dout[3]), .QN(n84) );
  DF3 Dout_reg_1_ ( .D(n103), .C(Clk), .Q(Dout[1]), .QN(n83) );
  DF3 Dout_reg_21_ ( .D(n65), .C(Clk), .Q(Dout[21]), .QN(n12) );
  DF3 Dout_reg_17_ ( .D(n69), .C(Clk), .Q(Dout[17]), .QN(n4) );
  DF3 Dout_reg_19_ ( .D(n67), .C(Clk), .Q(Dout[19]), .QN(n8) );
  DF3 Dout_reg_18_ ( .D(n68), .C(Clk), .Q(Dout[18]), .QN(n6) );
  DF3 Dout_reg_24_ ( .D(n62), .C(Clk), .Q(Dout[24]), .QN(n18) );
  DF3 Dout_reg_23_ ( .D(n63), .C(Clk), .Q(Dout[23]), .QN(n16) );
  DF3 Dout_reg_22_ ( .D(n64), .C(Clk), .Q(Dout[22]), .QN(n14) );
  DF3 Dout_reg_25_ ( .D(n61), .C(Clk), .Q(Dout[25]), .QN(n20) );
  OAI222 U3 ( .A(n82), .B(n360), .C(n362), .D(n368), .Q(n99) );
  OAI222 U4 ( .A(n76), .B(n360), .C(n361), .D(n370), .Q(n98) );
  OAI222 U5 ( .A(n77), .B(n360), .C(n109), .D(n371), .Q(n97) );
  OAI222 U6 ( .A(n78), .B(n360), .C(n362), .D(n377), .Q(n96) );
  OAI222 U7 ( .A(n79), .B(n360), .C(n361), .D(n378), .Q(n95) );
  OAI222 U8 ( .A(n80), .B(n360), .C(n109), .D(n376), .Q(n94) );
  OAI222 U9 ( .A(n81), .B(n360), .C(n362), .D(n375), .Q(n93) );
  OAI222 U10 ( .A(n71), .B(n360), .C(n361), .D(n379), .Q(n92) );
  OAI222 U11 ( .A(n72), .B(n360), .C(n109), .D(n374), .Q(n91) );
  OAI222 U12 ( .A(n73), .B(n360), .C(n362), .D(n373), .Q(n90) );
  OAI222 U13 ( .A(n74), .B(n360), .C(n361), .D(n372), .Q(n89) );
  OAI222 U14 ( .A(n87), .B(n360), .C(n109), .D(n381), .Q(n88) );
  OAI222 U15 ( .A(n4), .B(n360), .C(n362), .D(n394), .Q(n69) );
  OAI222 U16 ( .A(n6), .B(n360), .C(n361), .D(n384), .Q(n68) );
  OAI222 U17 ( .A(n8), .B(n360), .C(n109), .D(n385), .Q(n67) );
  OAI222 U18 ( .A(n10), .B(n360), .C(n362), .D(n380), .Q(n66) );
  OAI222 U19 ( .A(n12), .B(n360), .C(n361), .D(n395), .Q(n65) );
  OAI222 U20 ( .A(n14), .B(n360), .C(n109), .D(n387), .Q(n64) );
  OAI222 U21 ( .A(n16), .B(n360), .C(n362), .D(n386), .Q(n63) );
  OAI222 U22 ( .A(n18), .B(n360), .C(n361), .D(n383), .Q(n62) );
  OAI222 U23 ( .A(n20), .B(n360), .C(n109), .D(n390), .Q(n61) );
  OAI222 U24 ( .A(n22), .B(n360), .C(n362), .D(n393), .Q(n60) );
  OAI222 U25 ( .A(n24), .B(n360), .C(n361), .D(n389), .Q(n59) );
  OAI222 U26 ( .A(n26), .B(n360), .C(n109), .D(n391), .Q(n58) );
  OAI222 U27 ( .A(n28), .B(n360), .C(n362), .D(n388), .Q(n57) );
  OAI222 U28 ( .A(n30), .B(n360), .C(n361), .D(n382), .Q(n56) );
  OAI222 U29 ( .A(n32), .B(n360), .C(n392), .D(n109), .Q(n55) );
  OAI222 U30 ( .A(n86), .B(n360), .C(n362), .D(n364), .Q(n104) );
  OAI222 U31 ( .A(n83), .B(n360), .C(n361), .D(n365), .Q(n103) );
  OAI222 U32 ( .A(n75), .B(n360), .C(n109), .D(n367), .Q(n102) );
  OAI222 U33 ( .A(n84), .B(n360), .C(n362), .D(n366), .Q(n101) );
  OAI222 U34 ( .A(n85), .B(n360), .C(n361), .D(n369), .Q(n100) );
  DF1 Dout_reg_30_ ( .D(n56), .C(Clk), .Q(Dout[30]), .QN(n30) );
  DF1 Dout_reg_29_ ( .D(n57), .C(Clk), .Q(Dout[29]), .QN(n28) );
  DF1 Dout_reg_31_ ( .D(n55), .C(Clk), .Q(Dout[31]), .QN(n32) );
  DF3 Dout_reg_28_ ( .D(n58), .C(Clk), .Q(Dout[28]), .QN(n26) );
  DF3 Dout_reg_26_ ( .D(n60), .C(Clk), .Q(Dout[26]), .QN(n22) );
  DF3 Dout_reg_9_ ( .D(n95), .C(Clk), .Q(Dout[9]), .QN(n79) );
  DF3 Dout_reg_27_ ( .D(n59), .C(Clk), .Q(Dout[27]), .QN(n24) );
  DF3 Dout_reg_20_ ( .D(n66), .C(Clk), .Q(Dout[20]), .QN(n10) );
  INV4 U35 ( .A(Din[24]), .Q(n383) );
  INV3 U36 ( .A(Din[27]), .Q(n389) );
  INV3 U37 ( .A(Din[31]), .Q(n392) );
  INV3 U38 ( .A(Din[17]), .Q(n394) );
  INV3 U39 ( .A(Din[29]), .Q(n388) );
  INV3 U40 ( .A(Din[28]), .Q(n391) );
  INV3 U41 ( .A(Din[26]), .Q(n393) );
  INV3 U42 ( .A(Din[30]), .Q(n382) );
  INV4 U43 ( .A(Din[25]), .Q(n390) );
  INV3 U44 ( .A(Din[20]), .Q(n380) );
  INV2 U45 ( .A(Din[23]), .Q(n386) );
  INV2 U46 ( .A(Din[21]), .Q(n395) );
  INV2 U47 ( .A(Din[18]), .Q(n384) );
  INV2 U48 ( .A(Din[15]), .Q(n372) );
  INV2 U49 ( .A(Din[19]), .Q(n385) );
  INV2 U50 ( .A(Din[22]), .Q(n387) );
  INV2 U51 ( .A(Din[16]), .Q(n381) );
  INV2 U52 ( .A(Din[14]), .Q(n373) );
  INV2 U53 ( .A(Din[13]), .Q(n374) );
  NAND22 U54 ( .A(n363), .B(n360), .Q(n361) );
  NAND22 U55 ( .A(n363), .B(n360), .Q(n362) );
  NAND22 U56 ( .A(n363), .B(n360), .Q(n109) );
  INV3 U57 ( .A(Reset), .Q(n363) );
  INV3 U58 ( .A(n110), .Q(n360) );
  INV3 U59 ( .A(Din[12]), .Q(n379) );
  INV3 U60 ( .A(Din[8]), .Q(n377) );
  INV3 U61 ( .A(Din[11]), .Q(n375) );
  INV3 U62 ( .A(Din[10]), .Q(n376) );
  INV3 U63 ( .A(Din[9]), .Q(n378) );
  INV3 U64 ( .A(Din[7]), .Q(n371) );
  INV3 U65 ( .A(Din[3]), .Q(n366) );
  INV3 U66 ( .A(Din[4]), .Q(n369) );
  INV3 U67 ( .A(Din[5]), .Q(n368) );
  INV3 U68 ( .A(Din[6]), .Q(n370) );
  INV3 U69 ( .A(Din[2]), .Q(n367) );
  INV3 U70 ( .A(Din[1]), .Q(n365) );
  INV3 U71 ( .A(Din[0]), .Q(n364) );
  NOR20 U72 ( .A(Load), .B(Reset), .Q(n110) );
endmodule


module reg_8 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31,
         n34, n48, n50, n52, n54, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n56, n57, n58, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n107, n108, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393;

  DF3 Dout_reg_16_ ( .D(n74), .C(Clk), .Q(Dout[16]), .QN(n11) );
  DF3 Dout_reg_15_ ( .D(n75), .C(Clk), .Q(Dout[15]), .QN(n9) );
  DF3 Dout_reg_14_ ( .D(n76), .C(Clk), .Q(Dout[14]), .QN(n7) );
  DF3 Dout_reg_13_ ( .D(n77), .C(Clk), .Q(Dout[13]), .QN(n5) );
  DF3 Dout_reg_12_ ( .D(n88), .C(Clk), .Q(Dout[12]), .QN(n56) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n80) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n78) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n58) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n57) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n82) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n83) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n85) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n87) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n86) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n79) );
  DF3 Dout_reg_11_ ( .D(n89), .C(Clk), .Q(Dout[11]), .QN(n81) );
  DF3 Dout_reg_26_ ( .D(n64), .C(Clk), .Q(Dout[26]), .QN(n31) );
  DF3 Dout_reg_25_ ( .D(n65), .C(Clk), .Q(Dout[25]), .QN(n29) );
  OAI222 U3 ( .A(n86), .B(n358), .C(n360), .D(n393), .Q(n99) );
  OAI222 U4 ( .A(n85), .B(n358), .C(n359), .D(n390), .Q(n98) );
  OAI222 U5 ( .A(n84), .B(n358), .C(n107), .D(n391), .Q(n97) );
  OAI222 U6 ( .A(n83), .B(n358), .C(n360), .D(n388), .Q(n96) );
  OAI222 U7 ( .A(n82), .B(n358), .C(n359), .D(n389), .Q(n95) );
  OAI222 U8 ( .A(n57), .B(n358), .C(n107), .D(n386), .Q(n94) );
  OAI222 U9 ( .A(n58), .B(n358), .C(n360), .D(n387), .Q(n93) );
  OAI222 U10 ( .A(n78), .B(n358), .C(n359), .D(n385), .Q(n92) );
  OAI222 U11 ( .A(n79), .B(n358), .C(n107), .D(n384), .Q(n91) );
  OAI222 U12 ( .A(n80), .B(n358), .C(n360), .D(n383), .Q(n90) );
  OAI222 U13 ( .A(n81), .B(n358), .C(n359), .D(n380), .Q(n89) );
  OAI222 U14 ( .A(n56), .B(n358), .C(n107), .D(n382), .Q(n88) );
  OAI222 U15 ( .A(n5), .B(n358), .C(n360), .D(n381), .Q(n77) );
  OAI222 U16 ( .A(n7), .B(n358), .C(n359), .D(n379), .Q(n76) );
  OAI222 U17 ( .A(n9), .B(n358), .C(n107), .D(n378), .Q(n75) );
  OAI222 U18 ( .A(n11), .B(n358), .C(n360), .D(n377), .Q(n74) );
  OAI222 U19 ( .A(n13), .B(n358), .C(n359), .D(n376), .Q(n73) );
  OAI222 U20 ( .A(n15), .B(n358), .C(n107), .D(n375), .Q(n72) );
  OAI222 U21 ( .A(n17), .B(n358), .C(n360), .D(n374), .Q(n71) );
  OAI222 U22 ( .A(n19), .B(n358), .C(n359), .D(n373), .Q(n70) );
  OAI222 U23 ( .A(n21), .B(n358), .C(n372), .D(n107), .Q(n69) );
  OAI222 U24 ( .A(n23), .B(n358), .C(n360), .D(n371), .Q(n68) );
  OAI222 U25 ( .A(n25), .B(n358), .C(n359), .D(n370), .Q(n67) );
  OAI222 U26 ( .A(n27), .B(n358), .C(n107), .D(n369), .Q(n66) );
  OAI222 U27 ( .A(n29), .B(n358), .C(n368), .D(n360), .Q(n65) );
  OAI222 U28 ( .A(n31), .B(n358), .C(n367), .D(n359), .Q(n64) );
  OAI222 U29 ( .A(n34), .B(n358), .C(n366), .D(n107), .Q(n63) );
  OAI222 U30 ( .A(n48), .B(n358), .C(n365), .D(n360), .Q(n62) );
  OAI222 U31 ( .A(n50), .B(n358), .C(n364), .D(n359), .Q(n61) );
  OAI222 U32 ( .A(n52), .B(n358), .C(n107), .D(n363), .Q(n60) );
  OAI222 U33 ( .A(n54), .B(n358), .C(n362), .D(n360), .Q(n59) );
  OAI222 U34 ( .A(n87), .B(n358), .C(n359), .D(n392), .Q(n100) );
  DF1 Dout_reg_27_ ( .D(n63), .C(Clk), .Q(Dout[27]), .QN(n34) );
  DF1 Dout_reg_24_ ( .D(n66), .C(Clk), .Q(Dout[24]), .QN(n27) );
  DF1 Dout_reg_20_ ( .D(n70), .C(Clk), .Q(Dout[20]), .QN(n19) );
  DF1 Dout_reg_31_ ( .D(n59), .C(Clk), .Q(Dout[31]), .QN(n54) );
  DF1 Dout_reg_30_ ( .D(n60), .C(Clk), .Q(Dout[30]), .QN(n52) );
  DF1 Dout_reg_29_ ( .D(n61), .C(Clk), .Q(Dout[29]), .QN(n50) );
  DF3 Dout_reg_28_ ( .D(n62), .C(Clk), .Q(Dout[28]), .QN(n48) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n84) );
  DF3 Dout_reg_19_ ( .D(n71), .C(Clk), .Q(Dout[19]), .QN(n17) );
  DF3 Dout_reg_18_ ( .D(n72), .C(Clk), .Q(Dout[18]), .QN(n15) );
  DF3 Dout_reg_23_ ( .D(n67), .C(Clk), .Q(Dout[23]), .QN(n25) );
  DF3 Dout_reg_17_ ( .D(n73), .C(Clk), .Q(Dout[17]), .QN(n13) );
  DF3 Dout_reg_22_ ( .D(n68), .C(Clk), .Q(Dout[22]), .QN(n23) );
  DF3 Dout_reg_21_ ( .D(n69), .C(Clk), .Q(Dout[21]), .QN(n21) );
  INV4 U35 ( .A(Din[26]), .Q(n367) );
  INV4 U36 ( .A(Din[18]), .Q(n375) );
  INV4 U37 ( .A(Din[29]), .Q(n364) );
  INV4 U38 ( .A(Din[17]), .Q(n376) );
  INV3 U39 ( .A(Din[28]), .Q(n365) );
  INV3 U40 ( .A(Din[27]), .Q(n366) );
  INV4 U41 ( .A(Din[31]), .Q(n362) );
  INV4 U42 ( .A(Din[23]), .Q(n370) );
  INV3 U43 ( .A(Din[16]), .Q(n377) );
  INV3 U44 ( .A(Din[30]), .Q(n363) );
  CLKIN6 U45 ( .A(Din[21]), .Q(n372) );
  INV4 U46 ( .A(Din[25]), .Q(n368) );
  INV3 U47 ( .A(Din[22]), .Q(n371) );
  CLKIN3 U48 ( .A(Din[14]), .Q(n379) );
  INV2 U49 ( .A(Din[10]), .Q(n383) );
  INV2 U50 ( .A(Din[8]), .Q(n385) );
  INV2 U51 ( .A(Din[11]), .Q(n380) );
  CLKIN3 U52 ( .A(Din[12]), .Q(n382) );
  INV2 U53 ( .A(Din[9]), .Q(n384) );
  INV2 U54 ( .A(Din[24]), .Q(n369) );
  INV2 U55 ( .A(Din[20]), .Q(n373) );
  INV2 U56 ( .A(Din[19]), .Q(n374) );
  INV2 U57 ( .A(Din[13]), .Q(n381) );
  INV2 U58 ( .A(Din[15]), .Q(n378) );
  NAND22 U59 ( .A(n361), .B(n358), .Q(n359) );
  NAND22 U60 ( .A(n361), .B(n358), .Q(n360) );
  NAND22 U61 ( .A(n361), .B(n358), .Q(n107) );
  INV3 U62 ( .A(Reset), .Q(n361) );
  INV3 U63 ( .A(n108), .Q(n358) );
  INV3 U64 ( .A(Din[5]), .Q(n389) );
  INV3 U65 ( .A(Din[6]), .Q(n386) );
  INV3 U66 ( .A(Din[4]), .Q(n388) );
  INV3 U67 ( .A(Din[7]), .Q(n387) );
  INV3 U68 ( .A(Din[1]), .Q(n393) );
  INV3 U69 ( .A(Din[2]), .Q(n390) );
  INV3 U70 ( .A(Din[3]), .Q(n391) );
  INV3 U71 ( .A(Din[0]), .Q(n392) );
  NOR20 U72 ( .A(Load), .B(Reset), .Q(n108) );
endmodule


module adder_31_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n417, n418, n419,
         n420, n625, n626, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U59 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U219 ( .A(n787), .B(n197), .C(n419), .Q(n196) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U257 ( .A(n226), .B(n787), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n787), .B(n785), .C(n783), .Q(n232) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n271), .B(n275), .C(n272), .Q(n270) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U402 ( .A(n248), .B(n418), .C(n249), .Q(n420) );
  AOI212 U404 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U434 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U401 ( .A(n208), .B(n787), .C(n209), .Q(n207) );
  OAI212 U416 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U387 ( .A(n120), .B(n764), .C(n121), .Q(n119) );
  OAI212 U392 ( .A(n766), .B(n764), .C(n769), .Q(n164) );
  OAI212 U393 ( .A(n158), .B(n764), .C(n159), .Q(n157) );
  OAI212 U445 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U448 ( .A(n768), .B(n764), .C(n771), .Q(n108) );
  OAI212 U350 ( .A(n274), .B(n795), .C(n275), .Q(n273) );
  OAI212 U380 ( .A(n129), .B(n764), .C(n130), .Q(n128) );
  OAI212 U417 ( .A(n275), .B(n271), .C(n272), .Q(n417) );
  OAI212 U421 ( .A(n244), .B(n787), .C(n245), .Q(n243) );
  OAI212 U425 ( .A(n140), .B(n764), .C(n141), .Q(n139) );
  OAI212 U435 ( .A(n176), .B(n764), .C(n177), .Q(n175) );
  OAI212 U488 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U438 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U490 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U352 ( .A(n281), .B(n278), .C(n279), .Q(n625) );
  XNR22 U366 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NOR24 U409 ( .A(B[11]), .B(A[11]), .Q(n223) );
  OAI212 U413 ( .A(n91), .B(n764), .C(n92), .Q(n90) );
  OAI212 U422 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U429 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  XNR22 U437 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XNR22 U441 ( .A(n29), .B(n243), .Q(SUM[9]) );
  XNR22 U457 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U459 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U460 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U464 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U469 ( .A(n12), .B(n90), .Q(SUM[26]) );
  XNR22 U471 ( .A(n18), .B(n146), .Q(SUM[20]) );
  OAI212 U461 ( .A(n73), .B(n764), .C(n74), .Q(n72) );
  OAI212 U453 ( .A(n64), .B(n764), .C(n65), .Q(n63) );
  AOI212 U456 ( .A(n277), .B(n269), .C(n270), .Q(n418) );
  AOI212 U485 ( .A(n793), .B(n258), .C(n259), .Q(n257) );
  OAI212 U351 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  NOR24 U354 ( .A(B[4]), .B(A[4]), .Q(n265) );
  OAI212 U355 ( .A(n194), .B(n776), .C(n195), .Q(n191) );
  NOR24 U358 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR24 U370 ( .A(n185), .B(n194), .Q(n183) );
  NOR24 U412 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR24 U430 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR24 U431 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR24 U462 ( .A(n271), .B(n274), .Q(n269) );
  OAI212 U467 ( .A(n42), .B(n764), .C(n43), .Q(n41) );
  OAI212 U472 ( .A(n53), .B(n764), .C(n54), .Q(n52) );
  OAI212 U473 ( .A(n82), .B(n764), .C(n83), .Q(n81) );
  OAI212 U513 ( .A(n126), .B(n806), .C(n127), .Q(n123) );
  NOR23 U349 ( .A(B[7]), .B(A[7]), .Q(n252) );
  INV3 U353 ( .A(n230), .Q(n779) );
  OAI212 U356 ( .A(n102), .B(n764), .C(n103), .Q(n101) );
  NAND21 U357 ( .A(n111), .B(n809), .Q(n102) );
  XNR22 U359 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR22 U360 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NOR23 U361 ( .A(B[1]), .B(A[1]), .Q(n278) );
  XNR22 U362 ( .A(n225), .B(n27), .Q(SUM[11]) );
  NAND26 U363 ( .A(n135), .B(n115), .Q(n113) );
  AOI212 U364 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NOR22 U365 ( .A(n117), .B(n126), .Q(n115) );
  NAND24 U367 ( .A(n258), .B(n250), .Q(n248) );
  NOR22 U368 ( .A(n265), .B(n260), .Q(n258) );
  XNR22 U369 ( .A(n15), .B(n119), .Q(SUM[23]) );
  XOR22 U371 ( .A(n33), .B(n262), .Q(SUM[5]) );
  XNR22 U372 ( .A(n31), .B(n254), .Q(SUM[7]) );
  OAI211 U373 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  AOI212 U374 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  XNR22 U375 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XNR22 U376 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND21 U377 ( .A(n780), .B(n203), .Q(n197) );
  INV3 U378 ( .A(n219), .Q(n780) );
  XNR22 U379 ( .A(n20), .B(n164), .Q(SUM[18]) );
  XNR22 U381 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND22 U382 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NOR23 U383 ( .A(n219), .B(n181), .Q(n179) );
  NOR23 U384 ( .A(n252), .B(n255), .Q(n250) );
  NOR22 U385 ( .A(n99), .B(n106), .Q(n97) );
  NOR22 U386 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR22 U388 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR22 U389 ( .A(n173), .B(n176), .Q(n171) );
  INV3 U390 ( .A(n151), .Q(n767) );
  NOR23 U391 ( .A(n223), .B(n230), .Q(n221) );
  NAND22 U394 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND23 U395 ( .A(n171), .B(n153), .Q(n151) );
  NAND22 U396 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND22 U397 ( .A(n800), .B(n174), .Q(n21) );
  NOR21 U398 ( .A(n79), .B(n88), .Q(n77) );
  NOR21 U399 ( .A(n88), .B(n810), .Q(n84) );
  NOR23 U400 ( .A(n137), .B(n144), .Q(n135) );
  NOR23 U403 ( .A(B[10]), .B(A[10]), .Q(n230) );
  AOI211 U405 ( .A(n277), .B(n269), .C(n417), .Q(n268) );
  AOI211 U406 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR22 U407 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR22 U408 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR22 U410 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR22 U411 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NAND22 U414 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NOR22 U415 ( .A(B[21]), .B(A[21]), .Q(n137) );
  AOI211 U418 ( .A(n770), .B(n807), .C(n805), .Q(n141) );
  NOR23 U419 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NAND23 U420 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NOR22 U423 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND23 U424 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U426 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NOR22 U427 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND22 U428 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR23 U432 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NAND22 U433 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NOR22 U436 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR22 U439 ( .A(B[16]), .B(A[16]), .Q(n176) );
  XNR21 U440 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR21 U442 ( .A(n14), .B(n108), .Q(SUM[24]) );
  AOI211 U443 ( .A(n763), .B(n55), .C(n56), .Q(n54) );
  NOR21 U444 ( .A(n821), .B(n6), .Q(n55) );
  NOR21 U446 ( .A(n126), .B(n808), .Q(n122) );
  INV3 U447 ( .A(n135), .Q(n808) );
  AOI211 U449 ( .A(n781), .B(n190), .C(n191), .Q(n189) );
  AOI211 U450 ( .A(n625), .B(n269), .C(n270), .Q(n626) );
  INV2 U451 ( .A(n626), .Q(n793) );
  XOR21 U452 ( .A(n257), .B(n32), .Q(SUM[6]) );
  INV8 U454 ( .A(n420), .Q(n787) );
  INV2 U455 ( .A(n220), .Q(n781) );
  XOR22 U458 ( .A(n22), .B(n764), .Q(SUM[16]) );
  INV2 U463 ( .A(n152), .Q(n770) );
  NAND22 U465 ( .A(A[11]), .B(B[11]), .Q(n224) );
  AOI211 U466 ( .A(n809), .B(n763), .C(n812), .Q(n103) );
  NAND23 U468 ( .A(n239), .B(n221), .Q(n219) );
  NAND21 U470 ( .A(n239), .B(n779), .Q(n226) );
  NOR22 U474 ( .A(n241), .B(n244), .Q(n239) );
  NAND22 U475 ( .A(B[9]), .B(A[9]), .Q(n242) );
  NAND22 U476 ( .A(A[3]), .B(B[3]), .Q(n272) );
  AOI211 U477 ( .A(n781), .B(n777), .C(n778), .Q(n209) );
  AOI211 U478 ( .A(n781), .B(n203), .C(n204), .Q(n419) );
  OAI211 U479 ( .A(n188), .B(n787), .C(n189), .Q(n187) );
  AOI211 U480 ( .A(n763), .B(n811), .C(n814), .Q(n74) );
  INV6 U481 ( .A(n762), .Q(n763) );
  OAI211 U482 ( .A(n219), .B(n787), .C(n220), .Q(n214) );
  NAND22 U483 ( .A(A[23]), .B(B[23]), .Q(n118) );
  AOI211 U484 ( .A(n763), .B(n66), .C(n67), .Q(n65) );
  NAND22 U486 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NOR24 U487 ( .A(B[3]), .B(A[3]), .Q(n271) );
  OAI212 U489 ( .A(n151), .B(n764), .C(n152), .Q(n146) );
  NOR23 U491 ( .A(n155), .B(n162), .Q(n153) );
  NOR23 U492 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR24 U493 ( .A(n113), .B(n151), .Q(n111) );
  NAND22 U494 ( .A(n111), .B(n97), .Q(n91) );
  NAND22 U495 ( .A(n111), .B(n84), .Q(n82) );
  INV3 U496 ( .A(n111), .Q(n768) );
  NAND21 U497 ( .A(n111), .B(n55), .Q(n53) );
  NAND21 U498 ( .A(n111), .B(n44), .Q(n42) );
  NAND22 U499 ( .A(n767), .B(n135), .Q(n129) );
  INV1 U500 ( .A(n763), .Q(n771) );
  NAND22 U501 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NAND22 U502 ( .A(A[21]), .B(B[21]), .Q(n138) );
  CLKIN0 U503 ( .A(n173), .Q(n800) );
  NAND20 U504 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND21 U505 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND21 U506 ( .A(A[25]), .B(B[25]), .Q(n100) );
  INV1 U507 ( .A(n6), .Q(n811) );
  INV1 U508 ( .A(n5), .Q(n814) );
  CLKIN3 U509 ( .A(n60), .Q(n822) );
  INV0 U510 ( .A(n172), .Q(n769) );
  NAND21 U511 ( .A(n780), .B(n777), .Q(n208) );
  NAND21 U512 ( .A(n807), .B(n145), .Q(n18) );
  INV0 U514 ( .A(n212), .Q(n777) );
  XNR21 U515 ( .A(n34), .B(n793), .Q(SUM[4]) );
  INV0 U516 ( .A(n244), .Q(n784) );
  INV0 U517 ( .A(n204), .Q(n776) );
  AOI211 U518 ( .A(n793), .B(n790), .C(n791), .Q(n262) );
  INV3 U519 ( .A(n21), .Q(n761) );
  NAND22 U520 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR23 U521 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND22 U522 ( .A(B[1]), .B(A[1]), .Q(n279) );
  NAND22 U523 ( .A(n111), .B(n66), .Q(n64) );
  NAND21 U524 ( .A(n767), .B(n807), .Q(n140) );
  OAI210 U525 ( .A(n821), .B(n5), .C(n822), .Q(n56) );
  CLKIN0 U526 ( .A(n240), .Q(n783) );
  NAND21 U527 ( .A(n780), .B(n190), .Q(n188) );
  CLKIN3 U528 ( .A(n59), .Q(n821) );
  NAND20 U529 ( .A(n784), .B(n245), .Q(n30) );
  INV0 U530 ( .A(n61), .Q(n820) );
  INV0 U531 ( .A(n70), .Q(n827) );
  NOR23 U532 ( .A(n205), .B(n212), .Q(n203) );
  NAND20 U533 ( .A(n789), .B(n261), .Q(n33) );
  NAND20 U534 ( .A(n777), .B(n213), .Q(n26) );
  INV0 U535 ( .A(n265), .Q(n790) );
  AOI210 U536 ( .A(n60), .B(n818), .C(n817), .Q(n47) );
  NAND20 U537 ( .A(n792), .B(n275), .Q(n36) );
  INV0 U538 ( .A(n231), .Q(n782) );
  INV0 U539 ( .A(n98), .Q(n813) );
  OAI210 U540 ( .A(n88), .B(n813), .C(n89), .Q(n85) );
  NAND20 U541 ( .A(n790), .B(n266), .Q(n34) );
  INV0 U542 ( .A(n239), .Q(n785) );
  NAND20 U543 ( .A(n779), .B(n231), .Q(n28) );
  INV0 U544 ( .A(n79), .Q(n825) );
  NAND20 U545 ( .A(n825), .B(n80), .Q(n11) );
  INV0 U546 ( .A(n88), .Q(n819) );
  NAND20 U547 ( .A(n819), .B(n89), .Q(n12) );
  NAND22 U548 ( .A(n799), .B(n242), .Q(n29) );
  CLKIN0 U549 ( .A(n106), .Q(n809) );
  CLKIN0 U550 ( .A(n144), .Q(n807) );
  NAND20 U551 ( .A(n59), .B(n818), .Q(n46) );
  CLKIN0 U552 ( .A(n213), .Q(n778) );
  INV0 U553 ( .A(n271), .Q(n798) );
  NAND20 U554 ( .A(n798), .B(n272), .Q(n35) );
  CLKIN0 U555 ( .A(n97), .Q(n810) );
  INV0 U556 ( .A(n266), .Q(n791) );
  NOR24 U557 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR22 U558 ( .A(B[18]), .B(A[18]), .Q(n162) );
  INV2 U559 ( .A(n38), .Q(SUM[0]) );
  INV2 U560 ( .A(n280), .Q(n796) );
  NAND20 U561 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND21 U562 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND22 U563 ( .A(n111), .B(n811), .Q(n73) );
  NAND22 U564 ( .A(n97), .B(n77), .Q(n6) );
  NOR20 U565 ( .A(n46), .B(n6), .Q(n44) );
  AOI210 U566 ( .A(n770), .B(n135), .C(n136), .Q(n130) );
  NAND24 U567 ( .A(n203), .B(n183), .Q(n181) );
  INV1 U568 ( .A(n625), .Q(n795) );
  NAND22 U569 ( .A(n767), .B(n122), .Q(n120) );
  NAND20 U570 ( .A(n171), .B(n802), .Q(n158) );
  NAND22 U571 ( .A(n774), .B(n206), .Q(n25) );
  INV0 U572 ( .A(n205), .Q(n774) );
  NAND22 U573 ( .A(n804), .B(n118), .Q(n15) );
  INV3 U574 ( .A(n117), .Q(n804) );
  NAND22 U575 ( .A(n802), .B(n163), .Q(n20) );
  INV0 U576 ( .A(n171), .Q(n766) );
  NAND22 U577 ( .A(n816), .B(n138), .Q(n17) );
  INV3 U578 ( .A(n137), .Q(n816) );
  NAND22 U579 ( .A(n826), .B(n100), .Q(n13) );
  INV0 U580 ( .A(n99), .Q(n826) );
  NAND22 U581 ( .A(n815), .B(n224), .Q(n27) );
  INV0 U582 ( .A(n223), .Q(n815) );
  NAND22 U583 ( .A(n801), .B(n156), .Q(n19) );
  INV3 U584 ( .A(n155), .Q(n801) );
  NAND22 U585 ( .A(n824), .B(n127), .Q(n16) );
  INV3 U586 ( .A(n126), .Q(n824) );
  XOR22 U587 ( .A(n761), .B(n175), .Q(SUM[17]) );
  CLKIN0 U588 ( .A(n241), .Q(n799) );
  NAND22 U589 ( .A(n809), .B(n107), .Q(n14) );
  INV3 U590 ( .A(n107), .Q(n812) );
  NAND22 U591 ( .A(n788), .B(n256), .Q(n32) );
  INV0 U592 ( .A(n255), .Q(n788) );
  XOR21 U593 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U594 ( .A(n797), .B(n279), .Q(n37) );
  INV0 U595 ( .A(n278), .Q(n797) );
  XOR21 U596 ( .A(n787), .B(n30), .Q(SUM[8]) );
  NAND22 U597 ( .A(n765), .B(n177), .Q(n22) );
  INV0 U598 ( .A(n176), .Q(n765) );
  INV0 U599 ( .A(n260), .Q(n789) );
  XOR21 U600 ( .A(n36), .B(n795), .Q(SUM[2]) );
  INV0 U601 ( .A(n274), .Q(n792) );
  NAND22 U602 ( .A(n786), .B(n253), .Q(n31) );
  INV0 U603 ( .A(n252), .Q(n786) );
  NAND22 U604 ( .A(n772), .B(n186), .Q(n23) );
  INV0 U605 ( .A(n185), .Q(n772) );
  NAND22 U606 ( .A(n827), .B(n71), .Q(n10) );
  NAND22 U607 ( .A(n820), .B(n62), .Q(n9) );
  XNR21 U608 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND22 U609 ( .A(n818), .B(n51), .Q(n8) );
  INV3 U610 ( .A(n51), .Q(n817) );
  INV3 U611 ( .A(n163), .Q(n803) );
  XNR21 U612 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U613 ( .A(n773), .B(n195), .Q(n24) );
  INV0 U614 ( .A(n194), .Q(n773) );
  NOR21 U615 ( .A(n61), .B(n70), .Q(n59) );
  NOR21 U616 ( .A(n194), .B(n775), .Q(n190) );
  INV0 U617 ( .A(n203), .Q(n775) );
  NOR21 U618 ( .A(n70), .B(n6), .Q(n66) );
  AOI210 U619 ( .A(n770), .B(n122), .C(n123), .Q(n121) );
  INV0 U620 ( .A(n136), .Q(n806) );
  INV3 U621 ( .A(n145), .Q(n805) );
  INV3 U622 ( .A(n162), .Q(n802) );
  XNR21 U623 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U624 ( .A(n823), .B(n40), .Q(n7) );
  NAND22 U625 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR21 U626 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR21 U627 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND24 U628 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U629 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND21 U630 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND22 U631 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND22 U632 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND22 U633 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND22 U634 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV3 U635 ( .A(n50), .Q(n818) );
  NOR21 U636 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND20 U637 ( .A(n796), .B(n281), .Q(n38) );
  NOR20 U638 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U639 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U640 ( .A(n39), .Q(n823) );
  NOR21 U641 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV6 U642 ( .A(n112), .Q(n762) );
  AOI210 U643 ( .A(n172), .B(n802), .C(n803), .Q(n159) );
  AOI210 U644 ( .A(n240), .B(n779), .C(n782), .Q(n227) );
  CLKBU15 U645 ( .A(n178), .Q(n764) );
  AOI210 U646 ( .A(n763), .B(n44), .C(n45), .Q(n43) );
  AOI210 U647 ( .A(n763), .B(n84), .C(n85), .Q(n83) );
  AOI210 U648 ( .A(n763), .B(n97), .C(n98), .Q(n92) );
endmodule


module adder_31 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_31_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_30_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n420, n422,
         n430, n435, n436, n504, n576, n649, n786, n787, n788, n789, n790,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855;

  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n790), .C(n121), .Q(n119) );
  OAI212 U165 ( .A(n158), .B(n790), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n823), .B(n790), .C(n819), .Q(n164) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U233 ( .A(n208), .B(n795), .C(n209), .Q(n207) );
  OAI212 U257 ( .A(n226), .B(n795), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n810), .B(n795), .C(n808), .Q(n232) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U298 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n793), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U472 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U474 ( .A(n42), .B(n790), .C(n43), .Q(n41) );
  OAI212 U504 ( .A(n197), .B(n795), .C(n198), .Q(n196) );
  OAI212 U509 ( .A(n188), .B(n795), .C(n189), .Q(n187) );
  OAI212 U434 ( .A(n129), .B(n790), .C(n130), .Q(n128) );
  OAI212 U451 ( .A(n790), .B(n53), .C(n54), .Q(n52) );
  OAI212 U458 ( .A(n173), .B(n177), .C(n174), .Q(n172) );
  OAI212 U471 ( .A(n790), .B(n82), .C(n83), .Q(n81) );
  OAI212 U479 ( .A(n790), .B(n64), .C(n65), .Q(n63) );
  OAI212 U489 ( .A(n140), .B(n790), .C(n141), .Q(n139) );
  OAI212 U516 ( .A(n73), .B(n790), .C(n74), .Q(n72) );
  OAI212 U393 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  AOI212 U414 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U446 ( .A(n790), .B(n102), .C(n103), .Q(n101) );
  OAI212 U464 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U484 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U430 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U502 ( .A(n436), .B(n840), .C(n838), .Q(n56) );
  OAI212 U422 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U503 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U415 ( .A(n219), .B(n795), .C(n649), .Q(n214) );
  OAI212 U492 ( .A(n126), .B(n833), .C(n127), .Q(n123) );
  NAND24 U349 ( .A(n183), .B(n203), .Q(n181) );
  AOI211 U350 ( .A(n504), .B(n827), .C(n828), .Q(n159) );
  INV0 U351 ( .A(n171), .Q(n823) );
  CLKIN15 U352 ( .A(n788), .Q(n789) );
  NAND26 U353 ( .A(n420), .B(n80), .Q(n78) );
  NAND24 U354 ( .A(n845), .B(n850), .Q(n420) );
  NOR23 U355 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NAND26 U356 ( .A(n97), .B(n77), .Q(n6) );
  NOR23 U357 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR22 U358 ( .A(n212), .B(n205), .Q(n203) );
  INV3 U359 ( .A(n649), .Q(n805) );
  NAND23 U360 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NOR23 U361 ( .A(n117), .B(n126), .Q(n115) );
  NAND22 U362 ( .A(n430), .B(n224), .Q(n222) );
  NOR22 U363 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NAND22 U364 ( .A(n59), .B(n837), .Q(n46) );
  AOI211 U365 ( .A(n60), .B(n837), .C(n836), .Q(n47) );
  NOR22 U366 ( .A(n46), .B(n6), .Q(n44) );
  NOR23 U367 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR22 U368 ( .A(n173), .B(n176), .Q(n171) );
  NOR21 U369 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U370 ( .A(A[12]), .B(B[12]), .Q(n212) );
  AOI211 U371 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND22 U372 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND23 U373 ( .A(n576), .B(n786), .Q(n146) );
  NOR22 U374 ( .A(n840), .B(n6), .Q(n55) );
  NOR21 U375 ( .A(n194), .B(n816), .Q(n190) );
  XNR21 U376 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NOR24 U377 ( .A(A[21]), .B(B[21]), .Q(n137) );
  NAND22 U378 ( .A(A[21]), .B(B[21]), .Q(n138) );
  OAI212 U379 ( .A(n5), .B(n46), .C(n47), .Q(n45) );
  NAND22 U380 ( .A(n111), .B(n97), .Q(n91) );
  NAND26 U381 ( .A(n171), .B(n153), .Q(n151) );
  AOI212 U382 ( .A(n789), .B(n44), .C(n45), .Q(n43) );
  NAND21 U383 ( .A(n837), .B(n51), .Q(n8) );
  INV3 U384 ( .A(n820), .Q(n786) );
  CLKIN3 U385 ( .A(n152), .Q(n820) );
  AOI211 U386 ( .A(n805), .B(n190), .C(n191), .Q(n189) );
  INV6 U387 ( .A(n112), .Q(n788) );
  AOI212 U388 ( .A(n820), .B(n122), .C(n123), .Q(n121) );
  OAI212 U389 ( .A(n176), .B(n790), .C(n177), .Q(n175) );
  OAI210 U390 ( .A(n177), .B(n173), .C(n174), .Q(n504) );
  NAND20 U391 ( .A(n829), .B(n177), .Q(n22) );
  NAND22 U392 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND21 U394 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV2 U395 ( .A(n155), .Q(n826) );
  NAND20 U396 ( .A(n171), .B(n827), .Q(n158) );
  INV4 U397 ( .A(n151), .Q(n824) );
  NAND22 U398 ( .A(n122), .B(n824), .Q(n120) );
  BUF15 U399 ( .A(n178), .Q(n790) );
  NOR24 U400 ( .A(B[25]), .B(A[25]), .Q(n99) );
  CLKIN6 U401 ( .A(n79), .Q(n850) );
  NOR22 U402 ( .A(n88), .B(n854), .Q(n84) );
  INV1 U403 ( .A(n88), .Q(n842) );
  OAI211 U404 ( .A(n88), .B(n852), .C(n89), .Q(n85) );
  NOR23 U405 ( .A(n252), .B(n255), .Q(n250) );
  CLKIN3 U406 ( .A(n247), .Q(n795) );
  OAI211 U407 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  NAND21 U408 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NOR24 U409 ( .A(A[13]), .B(B[13]), .Q(n205) );
  CLKIN0 U410 ( .A(n204), .Q(n814) );
  INV0 U411 ( .A(n194), .Q(n817) );
  NAND20 U412 ( .A(n807), .B(n203), .Q(n197) );
  INV2 U413 ( .A(n203), .Q(n816) );
  NOR24 U416 ( .A(n61), .B(n70), .Q(n59) );
  AOI212 U417 ( .A(n789), .B(n66), .C(n67), .Q(n65) );
  AOI211 U418 ( .A(n820), .B(n834), .C(n832), .Q(n141) );
  AOI212 U419 ( .A(n789), .B(n84), .C(n85), .Q(n83) );
  NAND21 U420 ( .A(n853), .B(n107), .Q(n14) );
  OAI212 U421 ( .A(n107), .B(n99), .C(n100), .Q(n422) );
  XNR22 U423 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR22 U424 ( .A(n12), .B(n90), .Q(SUM[26]) );
  XNR22 U425 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XNR22 U426 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NAND21 U427 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV4 U428 ( .A(n59), .Q(n840) );
  OAI212 U429 ( .A(n436), .B(n70), .C(n71), .Q(n67) );
  XNR22 U431 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NOR24 U432 ( .A(A[22]), .B(B[22]), .Q(n126) );
  NOR24 U433 ( .A(n219), .B(n181), .Q(n179) );
  XOR21 U435 ( .A(n22), .B(n790), .Q(SUM[16]) );
  NAND26 U436 ( .A(n135), .B(n115), .Q(n113) );
  OAI212 U437 ( .A(n91), .B(n790), .C(n92), .Q(n90) );
  NOR24 U438 ( .A(n113), .B(n151), .Q(n111) );
  AOI212 U439 ( .A(n789), .B(n843), .C(n844), .Q(n74) );
  NOR24 U440 ( .A(n185), .B(n194), .Q(n183) );
  OAI210 U441 ( .A(n194), .B(n814), .C(n787), .Q(n191) );
  NOR24 U442 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR23 U443 ( .A(B[18]), .B(A[18]), .Q(n162) );
  XNR22 U444 ( .A(n7), .B(n41), .Q(SUM[31]) );
  CLKIN2 U445 ( .A(n60), .Q(n838) );
  INV0 U447 ( .A(n176), .Q(n829) );
  XNR22 U448 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR22 U449 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NOR24 U450 ( .A(A[26]), .B(B[26]), .Q(n88) );
  NOR24 U452 ( .A(n79), .B(n88), .Q(n77) );
  NAND21 U453 ( .A(A[15]), .B(B[15]), .Q(n186) );
  OAI212 U454 ( .A(n825), .B(n790), .C(n821), .Q(n108) );
  NOR22 U455 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR24 U456 ( .A(n99), .B(n106), .Q(n97) );
  NOR23 U457 ( .A(n155), .B(n162), .Q(n153) );
  AOI212 U459 ( .A(n435), .B(n115), .C(n116), .Q(n114) );
  NOR24 U460 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR24 U461 ( .A(n144), .B(n137), .Q(n135) );
  NAND22 U462 ( .A(A[22]), .B(B[22]), .Q(n127) );
  OAI212 U463 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND22 U465 ( .A(A[26]), .B(B[26]), .Q(n89) );
  AOI210 U466 ( .A(n805), .B(n203), .C(n204), .Q(n198) );
  AOI212 U467 ( .A(n789), .B(n853), .C(n851), .Q(n103) );
  NAND22 U468 ( .A(n111), .B(n853), .Q(n102) );
  INV1 U469 ( .A(n106), .Q(n853) );
  AOI212 U470 ( .A(n789), .B(n97), .C(n422), .Q(n92) );
  NAND21 U473 ( .A(B[23]), .B(A[23]), .Q(n118) );
  INV0 U475 ( .A(n145), .Q(n832) );
  OAI212 U476 ( .A(n137), .B(n145), .C(n138), .Q(n435) );
  NAND22 U477 ( .A(n111), .B(n843), .Q(n73) );
  INV3 U478 ( .A(n111), .Q(n825) );
  INV3 U480 ( .A(n6), .Q(n843) );
  INV1 U481 ( .A(n162), .Q(n827) );
  INV2 U482 ( .A(n97), .Q(n854) );
  INV1 U483 ( .A(n205), .Q(n815) );
  AOI211 U485 ( .A(n240), .B(n221), .C(n222), .Q(n649) );
  NAND22 U486 ( .A(A[27]), .B(B[27]), .Q(n80) );
  INV1 U487 ( .A(n144), .Q(n834) );
  NAND22 U488 ( .A(n111), .B(n44), .Q(n42) );
  NOR23 U490 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR24 U491 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR23 U493 ( .A(n241), .B(n244), .Q(n239) );
  OAI211 U494 ( .A(n244), .B(n795), .C(n245), .Q(n243) );
  INV0 U495 ( .A(n137), .Q(n849) );
  INV1 U496 ( .A(n789), .Q(n821) );
  NOR24 U497 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND22 U498 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND22 U499 ( .A(A[17]), .B(B[17]), .Q(n174) );
  CLKIN2 U500 ( .A(n135), .Q(n835) );
  AOI211 U501 ( .A(n820), .B(n135), .C(n136), .Q(n130) );
  XNR22 U505 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND21 U506 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NOR22 U507 ( .A(n70), .B(n6), .Q(n66) );
  NAND21 U508 ( .A(n847), .B(n71), .Q(n10) );
  NAND21 U510 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND22 U511 ( .A(B[25]), .B(A[25]), .Q(n100) );
  NAND24 U512 ( .A(B[16]), .B(A[16]), .Q(n177) );
  NAND21 U513 ( .A(n824), .B(n135), .Q(n129) );
  NAND21 U514 ( .A(n824), .B(n834), .Q(n140) );
  NAND21 U515 ( .A(B[10]), .B(A[10]), .Q(n231) );
  AOI212 U517 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  NOR23 U518 ( .A(n223), .B(n230), .Q(n221) );
  AOI212 U519 ( .A(n789), .B(n55), .C(n56), .Q(n54) );
  AOI212 U520 ( .A(n98), .B(n77), .C(n78), .Q(n436) );
  NAND21 U521 ( .A(n834), .B(n145), .Q(n18) );
  AOI212 U522 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  NAND24 U523 ( .A(n824), .B(n796), .Q(n576) );
  INV10 U524 ( .A(n790), .Q(n796) );
  NAND20 U525 ( .A(A[14]), .B(B[14]), .Q(n787) );
  INV3 U526 ( .A(n5), .Q(n844) );
  NOR22 U527 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR22 U528 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR22 U529 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NOR22 U530 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NAND20 U531 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NAND20 U532 ( .A(A[9]), .B(B[9]), .Q(n242) );
  INV0 U533 ( .A(n107), .Q(n851) );
  NAND21 U534 ( .A(A[12]), .B(B[12]), .Q(n213) );
  CLKIN3 U535 ( .A(n504), .Q(n819) );
  CLKIN0 U536 ( .A(n239), .Q(n810) );
  CLKIN0 U537 ( .A(n240), .Q(n808) );
  NAND22 U538 ( .A(n807), .B(n190), .Q(n188) );
  INV0 U539 ( .A(n163), .Q(n828) );
  INV2 U540 ( .A(n51), .Q(n836) );
  INV0 U541 ( .A(n212), .Q(n831) );
  NAND21 U542 ( .A(A[8]), .B(B[8]), .Q(n245) );
  INV2 U543 ( .A(n39), .Q(n848) );
  NAND21 U544 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND20 U545 ( .A(n239), .B(n812), .Q(n226) );
  NAND20 U546 ( .A(n258), .B(n250), .Q(n248) );
  INV0 U547 ( .A(n244), .Q(n809) );
  INV0 U548 ( .A(n252), .Q(n803) );
  NAND21 U549 ( .A(B[7]), .B(A[7]), .Q(n253) );
  NOR20 U550 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND20 U551 ( .A(n804), .B(n256), .Q(n32) );
  INV3 U552 ( .A(n219), .Q(n807) );
  AOI210 U553 ( .A(n240), .B(n812), .C(n813), .Q(n227) );
  NAND22 U554 ( .A(n239), .B(n221), .Q(n219) );
  AOI211 U555 ( .A(n794), .B(n258), .C(n259), .Q(n257) );
  INV3 U556 ( .A(n268), .Q(n794) );
  AOI211 U557 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U558 ( .A(n126), .B(n835), .Q(n122) );
  NAND22 U559 ( .A(n807), .B(n831), .Q(n208) );
  AOI210 U560 ( .A(n805), .B(n831), .C(n830), .Q(n209) );
  INV3 U561 ( .A(n213), .Q(n830) );
  INV3 U562 ( .A(n422), .Q(n852) );
  INV3 U563 ( .A(n136), .Q(n833) );
  NAND22 U564 ( .A(n813), .B(n806), .Q(n430) );
  INV3 U565 ( .A(n89), .Q(n845) );
  INV3 U566 ( .A(n230), .Q(n812) );
  INV3 U567 ( .A(n223), .Q(n806) );
  INV3 U568 ( .A(n173), .Q(n822) );
  INV3 U569 ( .A(n70), .Q(n847) );
  INV3 U570 ( .A(n99), .Q(n855) );
  INV3 U571 ( .A(n231), .Q(n813) );
  INV3 U572 ( .A(n61), .Q(n839) );
  INV3 U573 ( .A(n185), .Q(n818) );
  INV3 U574 ( .A(n117), .Q(n841) );
  NAND22 U575 ( .A(n803), .B(n253), .Q(n31) );
  INV3 U576 ( .A(n265), .Q(n800) );
  INV3 U577 ( .A(n255), .Q(n804) );
  NAND22 U578 ( .A(n798), .B(n272), .Q(n35) );
  INV3 U579 ( .A(n271), .Q(n798) );
  INV3 U580 ( .A(n241), .Q(n811) );
  NAND22 U581 ( .A(n802), .B(n261), .Q(n33) );
  INV3 U582 ( .A(n260), .Q(n802) );
  INV3 U583 ( .A(n274), .Q(n799) );
  INV3 U584 ( .A(n278), .Q(n797) );
  AOI211 U585 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U586 ( .A(n271), .B(n274), .Q(n269) );
  NOR21 U587 ( .A(n260), .B(n265), .Q(n258) );
  INV3 U588 ( .A(n277), .Q(n793) );
  INV3 U589 ( .A(n266), .Q(n801) );
  NOR21 U590 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND22 U591 ( .A(A[6]), .B(B[6]), .Q(n256) );
  INV3 U592 ( .A(n50), .Q(n837) );
  NOR21 U593 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NOR21 U594 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR21 U595 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U596 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U597 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U598 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U599 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U600 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U601 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U602 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND22 U603 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NOR21 U604 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U605 ( .A(n280), .Q(n792) );
  NOR21 U606 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U607 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U608 ( .A(n839), .B(n62), .Q(n9) );
  NAND20 U609 ( .A(n842), .B(n89), .Q(n12) );
  NAND20 U610 ( .A(n850), .B(n80), .Q(n11) );
  XNR21 U611 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U612 ( .A(n818), .B(n186), .Q(n23) );
  XNR21 U613 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U614 ( .A(n831), .B(n213), .Q(n26) );
  XNR21 U615 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U616 ( .A(n817), .B(n787), .Q(n24) );
  XOR21 U617 ( .A(n30), .B(n795), .Q(SUM[8]) );
  NAND20 U618 ( .A(n809), .B(n245), .Q(n30) );
  XNR21 U619 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U620 ( .A(n806), .B(n224), .Q(n27) );
  NAND22 U621 ( .A(n848), .B(n40), .Q(n7) );
  NAND20 U622 ( .A(n855), .B(n100), .Q(n13) );
  XNR21 U623 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U624 ( .A(n206), .B(n815), .Q(n25) );
  XNR21 U625 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U626 ( .A(n812), .B(n231), .Q(n28) );
  XNR21 U627 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U628 ( .A(n811), .B(n242), .Q(n29) );
  NAND20 U629 ( .A(n174), .B(n822), .Q(n21) );
  XNR21 U630 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND20 U631 ( .A(n846), .B(n127), .Q(n16) );
  XNR21 U632 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND20 U633 ( .A(n841), .B(n118), .Q(n15) );
  XNR21 U634 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND20 U635 ( .A(n827), .B(n163), .Q(n20) );
  XNR21 U636 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U637 ( .A(n826), .B(n156), .Q(n19) );
  XNR21 U638 ( .A(n17), .B(n139), .Q(SUM[21]) );
  NAND20 U639 ( .A(n138), .B(n849), .Q(n17) );
  XNR21 U640 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XNR21 U641 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XNR21 U642 ( .A(n34), .B(n794), .Q(SUM[4]) );
  NAND22 U643 ( .A(n800), .B(n266), .Q(n34) );
  XOR21 U644 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U645 ( .A(n794), .B(n800), .C(n801), .Q(n262) );
  XOR21 U646 ( .A(n32), .B(n257), .Q(SUM[6]) );
  XOR21 U647 ( .A(n36), .B(n793), .Q(SUM[2]) );
  NAND22 U648 ( .A(n799), .B(n275), .Q(n36) );
  XOR21 U649 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U650 ( .A(n797), .B(n279), .Q(n37) );
  INV3 U651 ( .A(n38), .Q(SUM[0]) );
  NAND22 U652 ( .A(n792), .B(n281), .Q(n38) );
  NAND22 U653 ( .A(n111), .B(n55), .Q(n53) );
  NAND22 U654 ( .A(n111), .B(n84), .Q(n82) );
  NAND22 U655 ( .A(n111), .B(n66), .Q(n64) );
  INV3 U656 ( .A(n126), .Q(n846) );
endmodule


module adder_30 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1, n3;

  adder_30_DW01_add_1 add_16 ( .A(A), .B({B[31:18], n3, B[16:0]}), .CI(n1), 
        .SUM(O) );
  BUF6 U1 ( .A(B[17]), .Q(n3) );
  LOGIC0 U2 ( .Q(n1) );
endmodule


module adder_29_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n423, n493,
         n494, n566, n567, n635, n636, n639, n641, n642, n780, n781, n782,
         n783, n784, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851;

  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U207 ( .A(n188), .B(n789), .C(n189), .Q(n187) );
  OAI212 U233 ( .A(n208), .B(n789), .C(n209), .Q(n207) );
  OAI212 U257 ( .A(n226), .B(n789), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n833), .B(n789), .C(n835), .Q(n232) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U298 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n787), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U406 ( .A(n120), .B(n784), .C(n121), .Q(n119) );
  OAI212 U407 ( .A(n140), .B(n784), .C(n141), .Q(n139) );
  OAI212 U420 ( .A(n849), .B(n784), .C(n847), .Q(n164) );
  OAI212 U421 ( .A(n158), .B(n784), .C(n159), .Q(n157) );
  OAI212 U435 ( .A(n129), .B(n784), .C(n130), .Q(n128) );
  OAI212 U409 ( .A(n42), .B(n784), .C(n43), .Q(n41) );
  OAI212 U413 ( .A(n102), .B(n784), .C(n103), .Q(n101) );
  OAI212 U440 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U404 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U484 ( .A(n126), .B(n818), .C(n127), .Q(n123) );
  OAI212 U492 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U375 ( .A(n82), .B(n784), .C(n83), .Q(n81) );
  AOI212 U418 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U422 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U472 ( .A(n176), .B(n784), .C(n177), .Q(n175) );
  OAI212 U400 ( .A(n219), .B(n789), .C(n494), .Q(n214) );
  AOI212 U437 ( .A(n240), .B(n221), .C(n222), .Q(n494) );
  OAI212 U457 ( .A(n73), .B(n784), .C(n74), .Q(n72) );
  OAI212 U462 ( .A(n64), .B(n784), .C(n65), .Q(n63) );
  OAI212 U469 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI212 U478 ( .A(n816), .B(n784), .C(n814), .Q(n108) );
  OAI212 U376 ( .A(n194), .B(n839), .C(n195), .Q(n191) );
  OAI212 U377 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  NOR24 U438 ( .A(A[13]), .B(B[13]), .Q(n205) );
  OAI212 U351 ( .A(n53), .B(n784), .C(n54), .Q(n52) );
  OAI212 U355 ( .A(n244), .B(n789), .C(n245), .Q(n243) );
  OAI212 U386 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U507 ( .A(n805), .B(n5), .C(n803), .Q(n56) );
  NOR21 U349 ( .A(n181), .B(n219), .Q(n179) );
  AOI211 U350 ( .A(n112), .B(n809), .C(n808), .Q(n74) );
  NOR23 U352 ( .A(n185), .B(n194), .Q(n183) );
  INV6 U353 ( .A(n247), .Q(n789) );
  NOR23 U354 ( .A(B[14]), .B(A[14]), .Q(n194) );
  OAI212 U356 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  XNR22 U357 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND22 U358 ( .A(n135), .B(n115), .Q(n113) );
  NOR22 U359 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NAND22 U360 ( .A(n10), .B(n72), .Q(n782) );
  NAND24 U361 ( .A(n780), .B(n781), .Q(n783) );
  NAND24 U362 ( .A(n782), .B(n783), .Q(SUM[28]) );
  INV6 U363 ( .A(n10), .Q(n780) );
  CLKIN6 U364 ( .A(n72), .Q(n781) );
  NOR20 U365 ( .A(B[2]), .B(A[2]), .Q(n274) );
  AOI212 U366 ( .A(n112), .B(n97), .C(n98), .Q(n92) );
  AOI211 U367 ( .A(n112), .B(n66), .C(n67), .Q(n65) );
  NAND26 U368 ( .A(n97), .B(n77), .Q(n6) );
  NOR23 U369 ( .A(n79), .B(n88), .Q(n77) );
  NOR22 U370 ( .A(n99), .B(n106), .Q(n97) );
  AOI211 U371 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  INV1 U372 ( .A(n230), .Q(n842) );
  NOR21 U373 ( .A(n117), .B(n126), .Q(n115) );
  INV3 U374 ( .A(n135), .Q(n820) );
  NOR23 U378 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR23 U379 ( .A(A[17]), .B(B[17]), .Q(n173) );
  INV3 U380 ( .A(n152), .Q(n824) );
  NOR21 U381 ( .A(n194), .B(n841), .Q(n190) );
  INV3 U382 ( .A(n231), .Q(n843) );
  INV3 U383 ( .A(n494), .Q(n836) );
  NOR21 U384 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR21 U385 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR21 U387 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR22 U388 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR22 U389 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR21 U390 ( .A(B[16]), .B(A[16]), .Q(n176) );
  XNR21 U391 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XNR21 U392 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XNR21 U393 ( .A(n26), .B(n214), .Q(SUM[12]) );
  AOI211 U394 ( .A(n112), .B(n831), .C(n830), .Q(n103) );
  AOI211 U395 ( .A(n112), .B(n55), .C(n56), .Q(n54) );
  AOI211 U396 ( .A(n836), .B(n190), .C(n191), .Q(n189) );
  NAND21 U397 ( .A(n842), .B(n231), .Q(n28) );
  CLKIN4 U398 ( .A(n157), .Q(n790) );
  OAI211 U399 ( .A(n197), .B(n789), .C(n198), .Q(n196) );
  OAI211 U401 ( .A(n245), .B(n241), .C(n242), .Q(n423) );
  INV2 U402 ( .A(n112), .Q(n814) );
  NOR23 U403 ( .A(n155), .B(n162), .Q(n153) );
  OAI212 U405 ( .A(n493), .B(n784), .C(n152), .Q(n146) );
  NOR20 U408 ( .A(B[1]), .B(A[1]), .Q(n278) );
  BUF15 U410 ( .A(n178), .Q(n784) );
  NAND22 U411 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NOR23 U412 ( .A(B[9]), .B(A[9]), .Q(n241) );
  XNR22 U414 ( .A(n27), .B(n225), .Q(SUM[11]) );
  OAI211 U415 ( .A(n91), .B(n784), .C(n92), .Q(n90) );
  NAND22 U416 ( .A(n832), .B(n245), .Q(n30) );
  NOR21 U417 ( .A(B[8]), .B(A[8]), .Q(n244) );
  OAI210 U419 ( .A(n213), .B(n205), .C(n206), .Q(n642) );
  OAI210 U423 ( .A(n213), .B(n205), .C(n206), .Q(n641) );
  NOR22 U424 ( .A(A[12]), .B(B[12]), .Q(n212) );
  XNR22 U425 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NAND22 U426 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND21 U427 ( .A(n819), .B(n138), .Q(n17) );
  OAI212 U428 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  INV1 U429 ( .A(n97), .Q(n812) );
  NAND22 U430 ( .A(n111), .B(n97), .Q(n91) );
  XNR22 U431 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NOR24 U432 ( .A(A[11]), .B(B[11]), .Q(n223) );
  NAND21 U433 ( .A(B[9]), .B(A[9]), .Q(n242) );
  NAND22 U434 ( .A(n826), .B(n135), .Q(n129) );
  NOR23 U436 ( .A(n137), .B(n144), .Q(n135) );
  XNR22 U439 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XNR22 U441 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NOR24 U442 ( .A(n223), .B(n230), .Q(n221) );
  CLKIN6 U443 ( .A(n223), .Q(n845) );
  INV1 U444 ( .A(n136), .Q(n818) );
  AOI211 U445 ( .A(n824), .B(n122), .C(n123), .Q(n121) );
  NOR22 U446 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR22 U447 ( .A(B[18]), .B(A[18]), .Q(n162) );
  XNR22 U448 ( .A(n9), .B(n63), .Q(SUM[29]) );
  AOI212 U449 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI211 U450 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NAND22 U451 ( .A(n111), .B(n55), .Q(n53) );
  NOR22 U452 ( .A(n805), .B(n6), .Q(n55) );
  NAND24 U453 ( .A(n635), .B(n636), .Q(SUM[19]) );
  NAND24 U454 ( .A(n566), .B(n567), .Q(SUM[17]) );
  NAND21 U455 ( .A(n21), .B(n175), .Q(n566) );
  NAND21 U456 ( .A(n826), .B(n122), .Q(n120) );
  NAND21 U458 ( .A(B[15]), .B(A[15]), .Q(n186) );
  XNR22 U459 ( .A(n20), .B(n164), .Q(SUM[18]) );
  CLKIN1 U460 ( .A(n203), .Q(n841) );
  XNR22 U461 ( .A(n23), .B(n187), .Q(SUM[15]) );
  XNR22 U463 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND22 U464 ( .A(A[13]), .B(B[13]), .Q(n206) );
  XNR22 U465 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND24 U466 ( .A(n639), .B(n224), .Q(n222) );
  NAND21 U467 ( .A(B[11]), .B(A[11]), .Q(n224) );
  INV3 U468 ( .A(n6), .Q(n809) );
  INV0 U470 ( .A(n185), .Q(n829) );
  NAND21 U471 ( .A(A[17]), .B(B[17]), .Q(n174) );
  XOR21 U473 ( .A(n22), .B(n784), .Q(SUM[16]) );
  NOR24 U474 ( .A(n113), .B(n151), .Q(n111) );
  NAND21 U475 ( .A(n111), .B(n831), .Q(n102) );
  NAND22 U476 ( .A(n111), .B(n66), .Q(n64) );
  NAND22 U477 ( .A(n111), .B(n84), .Q(n82) );
  CLKIN3 U479 ( .A(n111), .Q(n816) );
  NAND21 U480 ( .A(n111), .B(n809), .Q(n73) );
  NAND21 U481 ( .A(n111), .B(n44), .Q(n42) );
  XNR22 U482 ( .A(n17), .B(n139), .Q(SUM[21]) );
  INV1 U483 ( .A(n241), .Q(n837) );
  NOR20 U485 ( .A(n241), .B(n244), .Q(n239) );
  XNR22 U486 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND21 U487 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR22 U488 ( .A(B[20]), .B(A[20]), .Q(n144) );
  OAI210 U489 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  CLKIN1 U490 ( .A(n19), .Q(n823) );
  NAND21 U491 ( .A(n19), .B(n157), .Q(n635) );
  INV3 U493 ( .A(n423), .Q(n835) );
  NAND21 U494 ( .A(n810), .B(n89), .Q(n12) );
  NAND21 U495 ( .A(n806), .B(n71), .Q(n10) );
  NAND20 U496 ( .A(n831), .B(n107), .Q(n14) );
  INV0 U497 ( .A(n126), .Q(n817) );
  INV2 U498 ( .A(n244), .Q(n832) );
  NOR21 U499 ( .A(n61), .B(n70), .Q(n59) );
  NAND20 U500 ( .A(n239), .B(n842), .Q(n226) );
  NAND22 U501 ( .A(n799), .B(n253), .Q(n31) );
  INV2 U502 ( .A(n252), .Q(n799) );
  NAND20 U503 ( .A(n815), .B(n118), .Q(n15) );
  NAND21 U504 ( .A(A[18]), .B(B[18]), .Q(n163) );
  INV3 U505 ( .A(n5), .Q(n808) );
  NAND20 U506 ( .A(n834), .B(n203), .Q(n197) );
  NAND20 U508 ( .A(n834), .B(n840), .Q(n208) );
  NOR22 U509 ( .A(n173), .B(n176), .Q(n171) );
  INV0 U510 ( .A(n176), .Q(n851) );
  NAND20 U511 ( .A(n821), .B(n145), .Q(n18) );
  INV0 U512 ( .A(n213), .Q(n838) );
  NAND20 U513 ( .A(n171), .B(n828), .Q(n158) );
  INV1 U514 ( .A(n98), .Q(n813) );
  OAI210 U515 ( .A(n88), .B(n813), .C(n89), .Q(n85) );
  INV0 U516 ( .A(n99), .Q(n811) );
  INV0 U517 ( .A(n88), .Q(n810) );
  INV0 U518 ( .A(n70), .Q(n806) );
  NAND20 U519 ( .A(n817), .B(n127), .Q(n16) );
  CLKIN0 U520 ( .A(n172), .Q(n847) );
  NAND20 U521 ( .A(n828), .B(n163), .Q(n20) );
  INV0 U522 ( .A(n117), .Q(n815) );
  NAND20 U523 ( .A(n844), .B(n195), .Q(n24) );
  NAND20 U524 ( .A(n837), .B(n242), .Q(n29) );
  NAND20 U525 ( .A(n845), .B(n224), .Q(n27) );
  INV0 U526 ( .A(n155), .Q(n825) );
  NAND20 U527 ( .A(n59), .B(n802), .Q(n46) );
  CLKIN0 U528 ( .A(n106), .Q(n831) );
  NAND20 U529 ( .A(n840), .B(n213), .Q(n26) );
  NAND20 U530 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NOR22 U531 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND20 U532 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND20 U533 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NOR20 U534 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR20 U535 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND20 U536 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND21 U537 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND20 U538 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U539 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND20 U540 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NOR20 U541 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND20 U542 ( .A(A[4]), .B(B[4]), .Q(n266) );
  INV3 U543 ( .A(n493), .Q(n826) );
  INV3 U544 ( .A(n219), .Q(n834) );
  NAND22 U545 ( .A(n171), .B(n153), .Q(n151) );
  NOR20 U546 ( .A(n6), .B(n46), .Q(n44) );
  INV3 U547 ( .A(n60), .Q(n803) );
  AOI210 U548 ( .A(n824), .B(n135), .C(n136), .Q(n130) );
  AOI211 U549 ( .A(n423), .B(n842), .C(n843), .Q(n227) );
  NAND22 U550 ( .A(n171), .B(n153), .Q(n493) );
  NAND22 U551 ( .A(n846), .B(n791), .Q(n567) );
  INV3 U552 ( .A(n21), .Q(n846) );
  NAND22 U553 ( .A(n823), .B(n790), .Q(n636) );
  INV3 U554 ( .A(n175), .Q(n791) );
  NAND22 U555 ( .A(n203), .B(n183), .Q(n181) );
  NAND22 U556 ( .A(n826), .B(n821), .Q(n140) );
  INV3 U557 ( .A(n59), .Q(n805) );
  INV3 U558 ( .A(n171), .Q(n849) );
  AOI211 U559 ( .A(n788), .B(n258), .C(n259), .Q(n257) );
  NAND22 U560 ( .A(n239), .B(n221), .Q(n219) );
  INV3 U561 ( .A(n268), .Q(n788) );
  INV3 U562 ( .A(n277), .Q(n787) );
  NAND22 U563 ( .A(n834), .B(n190), .Q(n188) );
  NAND22 U564 ( .A(n851), .B(n177), .Q(n22) );
  AOI210 U565 ( .A(n172), .B(n828), .C(n827), .Q(n159) );
  INV3 U566 ( .A(n163), .Q(n827) );
  NAND22 U567 ( .A(n811), .B(n100), .Q(n13) );
  INV3 U568 ( .A(n239), .Q(n833) );
  XNR21 U569 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NOR23 U570 ( .A(n205), .B(n212), .Q(n203) );
  XOR21 U571 ( .A(n30), .B(n789), .Q(SUM[8]) );
  XOR21 U572 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND22 U573 ( .A(n798), .B(n256), .Q(n32) );
  INV3 U574 ( .A(n255), .Q(n798) );
  INV3 U575 ( .A(n137), .Q(n819) );
  XNR21 U576 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND22 U577 ( .A(n850), .B(n206), .Q(n25) );
  CLKIN0 U578 ( .A(n205), .Q(n850) );
  XNR21 U579 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND22 U580 ( .A(n807), .B(n80), .Q(n11) );
  INV3 U581 ( .A(n79), .Q(n807) );
  NAND22 U582 ( .A(n804), .B(n62), .Q(n9) );
  INV3 U583 ( .A(n61), .Q(n804) );
  NAND22 U584 ( .A(n802), .B(n51), .Q(n8) );
  NAND22 U585 ( .A(n829), .B(n186), .Q(n23) );
  NOR21 U586 ( .A(n126), .B(n820), .Q(n122) );
  AOI211 U587 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR21 U588 ( .A(n88), .B(n812), .Q(n84) );
  NOR21 U589 ( .A(n70), .B(n6), .Q(n66) );
  INV0 U590 ( .A(n194), .Q(n844) );
  INV3 U591 ( .A(n107), .Q(n830) );
  AOI210 U592 ( .A(n112), .B(n44), .C(n45), .Q(n43) );
  AOI211 U593 ( .A(n60), .B(n802), .C(n801), .Q(n47) );
  INV3 U594 ( .A(n51), .Q(n801) );
  AOI210 U595 ( .A(n836), .B(n203), .C(n642), .Q(n198) );
  NAND22 U596 ( .A(n848), .B(n174), .Q(n21) );
  INV3 U597 ( .A(n173), .Q(n848) );
  INV3 U598 ( .A(n641), .Q(n839) );
  AOI211 U599 ( .A(n824), .B(n821), .C(n822), .Q(n141) );
  INV3 U600 ( .A(n145), .Q(n822) );
  AOI211 U601 ( .A(n836), .B(n840), .C(n838), .Q(n209) );
  NAND22 U602 ( .A(n825), .B(n156), .Q(n19) );
  INV3 U603 ( .A(n144), .Q(n821) );
  NAND22 U604 ( .A(n843), .B(n845), .Q(n639) );
  INV3 U605 ( .A(n162), .Q(n828) );
  INV3 U606 ( .A(n212), .Q(n840) );
  XOR21 U607 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U608 ( .A(n788), .B(n796), .C(n795), .Q(n262) );
  NAND22 U609 ( .A(n797), .B(n261), .Q(n33) );
  INV3 U610 ( .A(n266), .Q(n795) );
  XNR21 U611 ( .A(n34), .B(n788), .Q(SUM[4]) );
  NAND22 U612 ( .A(n796), .B(n266), .Q(n34) );
  INV3 U613 ( .A(n260), .Q(n797) );
  XOR21 U614 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U615 ( .A(n792), .B(n279), .Q(n37) );
  INV3 U616 ( .A(n278), .Q(n792) );
  INV3 U617 ( .A(n265), .Q(n796) );
  XOR21 U618 ( .A(n36), .B(n787), .Q(SUM[2]) );
  NAND22 U619 ( .A(n793), .B(n275), .Q(n36) );
  INV3 U620 ( .A(n274), .Q(n793) );
  XNR21 U621 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U622 ( .A(n794), .B(n272), .Q(n35) );
  INV3 U623 ( .A(n271), .Q(n794) );
  AOI211 U624 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U625 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U626 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U627 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U628 ( .A(n252), .B(n255), .Q(n250) );
  NOR21 U629 ( .A(n260), .B(n265), .Q(n258) );
  NAND22 U630 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND22 U631 ( .A(B[10]), .B(A[10]), .Q(n231) );
  NOR21 U632 ( .A(B[28]), .B(A[28]), .Q(n70) );
  XNR21 U633 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U634 ( .A(n800), .B(n40), .Q(n7) );
  NAND22 U635 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND22 U636 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NOR21 U637 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR21 U638 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND22 U639 ( .A(B[8]), .B(A[8]), .Q(n245) );
  NAND21 U640 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND21 U641 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NOR20 U642 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR20 U643 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV3 U644 ( .A(n50), .Q(n802) );
  INV3 U645 ( .A(n39), .Q(n800) );
  NOR21 U646 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U647 ( .A(n38), .Q(SUM[0]) );
  NAND22 U648 ( .A(n786), .B(n281), .Q(n38) );
  INV3 U649 ( .A(n280), .Q(n786) );
  NOR20 U650 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U651 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U652 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND20 U653 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U654 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U655 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND20 U656 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND20 U657 ( .A(A[3]), .B(B[3]), .Q(n272) );
  AOI211 U658 ( .A(n112), .B(n84), .C(n85), .Q(n83) );
  NOR21 U659 ( .A(B[5]), .B(A[5]), .Q(n260) );
endmodule


module adder_29 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_29_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_28_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n43, n44, n47, n48,
         n49, n50, n51, n52, n55, n56, n57, n58, n59, n60, n63, n64, n65, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n82, n83, n84,
         n85, n86, n87, n92, n93, n94, n95, n96, n99, n100, n101, n102, n103,
         n109, n110, n111, n112, n113, n114, n117, n118, n119, n122, n123,
         n128, n129, n130, n131, n132, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n150, n151, n152,
         n153, n154, n155, n160, n161, n162, n163, n164, n167, n168, n169,
         n170, n171, n176, n177, n178, n179, n180, n181, n182, n185, n186,
         n187, n190, n191, n196, n197, n198, n199, n200, n202, n203, n204,
         n205, n206, n207, n208, n209, n211, n212, n215, n216, n217, n218,
         n223, n224, n225, n228, n229, n231, n232, n233, n234, n235, n236,
         n237, n238, n240, n241, n242, n245, n246, n247, n250, n251, n253,
         n254, n255, n256, n257, n258, n259, n260, n262, n263, n264, n265,
         n266, n403, n404, n483, n484, n554, n555, n773, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843;

  OAI212 U48 ( .A(n68), .B(n103), .C(n69), .Q(n2) );
  AOI212 U100 ( .A(n123), .B(n811), .C(n109), .Q(n103) );
  OAI212 U108 ( .A(n113), .B(n773), .C(n114), .Q(n112) );
  OAI212 U140 ( .A(n136), .B(n171), .C(n137), .Q(n135) );
  OAI212 U176 ( .A(n163), .B(n780), .C(n164), .Q(n162) );
  AOI212 U192 ( .A(n191), .B(n176), .C(n177), .Q(n171) );
  OAI212 U200 ( .A(n181), .B(n780), .C(n182), .Q(n180) );
  OAI212 U210 ( .A(n829), .B(n780), .C(n827), .Q(n187) );
  OAI212 U231 ( .A(n203), .B(n231), .C(n204), .Q(n202) );
  OAI212 U280 ( .A(n237), .B(n778), .C(n238), .Q(n236) );
  OAI212 U287 ( .A(n241), .B(n253), .C(n242), .Q(n240) );
  OAI212 U308 ( .A(n260), .B(n256), .C(n257), .Q(n255) );
  OAI212 U314 ( .A(n259), .B(n776), .C(n260), .Q(n258) );
  OAI212 U321 ( .A(n266), .B(n263), .C(n264), .Q(n262) );
  OAI212 U395 ( .A(n816), .B(n773), .C(n817), .Q(n119) );
  OAI212 U396 ( .A(n84), .B(n773), .C(n85), .Q(n83) );
  OAI212 U402 ( .A(n802), .B(n773), .C(n801), .Q(n65) );
  OAI212 U420 ( .A(n59), .B(n773), .C(n60), .Q(n58) );
  OAI212 U457 ( .A(n39), .B(n773), .C(n40), .Q(n38) );
  OAI212 U339 ( .A(n132), .B(n128), .C(n129), .Q(n123) );
  OAI212 U449 ( .A(n200), .B(n196), .C(n197), .Q(n191) );
  AOI212 U488 ( .A(n232), .B(n240), .C(n233), .Q(n231) );
  OAI212 U425 ( .A(n131), .B(n773), .C(n132), .Q(n130) );
  AOI212 U472 ( .A(n202), .B(n134), .C(n135), .Q(n1) );
  OAI212 U458 ( .A(n229), .B(n223), .C(n224), .Q(n218) );
  OAI212 U473 ( .A(n64), .B(n56), .C(n57), .Q(n55) );
  OAI212 U370 ( .A(n95), .B(n773), .C(n96), .Q(n94) );
  OAI212 U386 ( .A(n168), .B(n160), .C(n161), .Q(n155) );
  OAI212 U403 ( .A(n102), .B(n773), .C(n103), .Q(n101) );
  OAI212 U421 ( .A(n75), .B(n773), .C(n76), .Q(n74) );
  OAI212 U466 ( .A(n82), .B(n72), .C(n73), .Q(n71) );
  INV2 U334 ( .A(n171), .Q(n826) );
  CLKIN3 U335 ( .A(n212), .Q(n841) );
  NAND21 U336 ( .A(n810), .B(n86), .Q(n84) );
  NOR24 U337 ( .A(n160), .B(n167), .Q(n154) );
  XNR22 U338 ( .A(n6), .B(n58), .Q(SUM[29]) );
  XOR22 U340 ( .A(n15), .B(n773), .Q(SUM[20]) );
  NAND22 U341 ( .A(n810), .B(n77), .Q(n75) );
  NOR22 U342 ( .A(n79), .B(n805), .Q(n77) );
  CLKIN2 U343 ( .A(n86), .Q(n805) );
  NOR22 U344 ( .A(n128), .B(n131), .Q(n122) );
  NOR22 U345 ( .A(B[21]), .B(A[21]), .Q(n128) );
  NAND24 U346 ( .A(n190), .B(n176), .Q(n170) );
  NOR22 U347 ( .A(n196), .B(n199), .Q(n190) );
  NOR21 U348 ( .A(n56), .B(n63), .Q(n52) );
  NAND23 U349 ( .A(n122), .B(n811), .Q(n102) );
  NOR21 U350 ( .A(B[23]), .B(A[23]), .Q(n110) );
  NOR22 U351 ( .A(B[17]), .B(A[17]), .Q(n160) );
  NOR22 U352 ( .A(B[14]), .B(A[14]), .Q(n185) );
  INV3 U353 ( .A(n74), .Q(n782) );
  AOI211 U354 ( .A(n809), .B(n86), .C(n87), .Q(n85) );
  NOR21 U355 ( .A(B[25]), .B(A[25]), .Q(n92) );
  AOI211 U356 ( .A(n826), .B(n822), .C(n820), .Q(n164) );
  NOR22 U357 ( .A(n223), .B(n228), .Q(n217) );
  INV6 U358 ( .A(n202), .Q(n780) );
  XNR21 U359 ( .A(n7), .B(n65), .Q(SUM[28]) );
  XNR21 U360 ( .A(n5), .B(n49), .Q(SUM[30]) );
  NAND22 U361 ( .A(n837), .B(n229), .Q(n27) );
  NOR22 U362 ( .A(B[11]), .B(A[11]), .Q(n207) );
  NOR22 U363 ( .A(n212), .B(n207), .Q(n205) );
  NAND21 U364 ( .A(n818), .B(n141), .Q(n16) );
  NOR22 U365 ( .A(A[10]), .B(B[10]), .Q(n212) );
  OAI211 U366 ( .A(n50), .B(n773), .C(n51), .Q(n49) );
  NAND22 U367 ( .A(A[26]), .B(B[26]), .Q(n82) );
  INV1 U368 ( .A(n218), .Q(n836) );
  NAND20 U369 ( .A(n842), .B(n224), .Q(n26) );
  NOR22 U371 ( .A(B[16]), .B(A[16]), .Q(n167) );
  NAND21 U372 ( .A(n843), .B(n197), .Q(n22) );
  NOR21 U373 ( .A(B[22]), .B(A[22]), .Q(n117) );
  XNR22 U374 ( .A(n11), .B(n101), .Q(SUM[24]) );
  XOR22 U375 ( .A(n23), .B(n780), .Q(SUM[12]) );
  NAND22 U376 ( .A(n8), .B(n74), .Q(n554) );
  NAND22 U377 ( .A(A[24]), .B(B[24]), .Q(n100) );
  NAND21 U378 ( .A(A[15]), .B(B[15]), .Q(n179) );
  XOR22 U379 ( .A(n24), .B(n209), .Q(SUM[11]) );
  AOI210 U380 ( .A(n826), .B(n154), .C(n155), .Q(n153) );
  CLKIN3 U381 ( .A(n168), .Q(n820) );
  AOI212 U382 ( .A(n155), .B(n138), .C(n139), .Q(n137) );
  NOR20 U383 ( .A(A[7]), .B(B[7]), .Q(n234) );
  INV1 U384 ( .A(n154), .Q(n823) );
  NAND21 U385 ( .A(B[9]), .B(A[9]), .Q(n224) );
  NAND22 U387 ( .A(A[14]), .B(B[14]), .Q(n186) );
  AOI212 U388 ( .A(n205), .B(n218), .C(n206), .Q(n204) );
  NOR23 U389 ( .A(B[9]), .B(A[9]), .Q(n223) );
  NAND24 U390 ( .A(n799), .B(n782), .Q(n555) );
  NAND28 U391 ( .A(n554), .B(n555), .Q(SUM[27]) );
  XNR22 U392 ( .A(n17), .B(n151), .Q(SUM[18]) );
  NOR21 U393 ( .A(B[29]), .B(A[29]), .Q(n56) );
  XNR22 U394 ( .A(n20), .B(n180), .Q(SUM[15]) );
  BUF15 U397 ( .A(n1), .Q(n773) );
  OAI212 U398 ( .A(n199), .B(n780), .C(n200), .Q(n198) );
  NAND22 U399 ( .A(A[10]), .B(B[10]), .Q(n215) );
  INV2 U400 ( .A(n102), .Q(n810) );
  INV6 U401 ( .A(n404), .Q(n811) );
  XNR22 U404 ( .A(n22), .B(n198), .Q(SUM[13]) );
  OAI211 U405 ( .A(n212), .B(n836), .C(n215), .Q(n211) );
  XNR22 U406 ( .A(n9), .B(n83), .Q(SUM[26]) );
  OAI212 U407 ( .A(n100), .B(n92), .C(n93), .Q(n87) );
  OAI212 U408 ( .A(n207), .B(n215), .C(n208), .Q(n206) );
  NOR24 U409 ( .A(B[13]), .B(A[13]), .Q(n196) );
  OAI211 U410 ( .A(n152), .B(n780), .C(n153), .Q(n151) );
  AOI211 U411 ( .A(n779), .B(n217), .C(n218), .Q(n216) );
  AOI212 U412 ( .A(n779), .B(n837), .C(n835), .Q(n225) );
  AOI212 U413 ( .A(n779), .B(n838), .C(n211), .Q(n209) );
  XNR21 U414 ( .A(n27), .B(n779), .Q(SUM[8]) );
  INV2 U415 ( .A(n231), .Q(n779) );
  XOR22 U416 ( .A(n25), .B(n216), .Q(SUM[10]) );
  OAI212 U417 ( .A(n186), .B(n178), .C(n179), .Q(n177) );
  NAND21 U418 ( .A(B[17]), .B(A[17]), .Q(n161) );
  INV1 U419 ( .A(n155), .Q(n821) );
  NAND21 U422 ( .A(n832), .B(n186), .Q(n21) );
  OAI211 U423 ( .A(n170), .B(n780), .C(n171), .Q(n169) );
  CLKIN3 U424 ( .A(n186), .Q(n831) );
  INV1 U426 ( .A(n196), .Q(n843) );
  NOR22 U427 ( .A(n72), .B(n79), .Q(n70) );
  OAI210 U428 ( .A(n79), .B(n806), .C(n82), .Q(n78) );
  INV1 U429 ( .A(n79), .Q(n803) );
  NAND24 U430 ( .A(n86), .B(n70), .Q(n68) );
  NOR22 U431 ( .A(B[8]), .B(A[8]), .Q(n228) );
  NAND21 U432 ( .A(n825), .B(n822), .Q(n163) );
  NAND20 U433 ( .A(n822), .B(n168), .Q(n19) );
  INV1 U434 ( .A(n167), .Q(n822) );
  NAND22 U435 ( .A(A[12]), .B(B[12]), .Q(n200) );
  XNR22 U436 ( .A(n12), .B(n112), .Q(SUM[23]) );
  NAND21 U437 ( .A(A[11]), .B(B[11]), .Q(n208) );
  NAND22 U438 ( .A(A[8]), .B(B[8]), .Q(n229) );
  INV0 U439 ( .A(n100), .Q(n807) );
  AOI212 U440 ( .A(n87), .B(n70), .C(n71), .Q(n69) );
  XNR22 U441 ( .A(n21), .B(n187), .Q(SUM[14]) );
  XNR22 U442 ( .A(n16), .B(n142), .Q(SUM[19]) );
  OAI211 U443 ( .A(n143), .B(n780), .C(n144), .Q(n142) );
  NAND22 U444 ( .A(n3), .B(n52), .Q(n50) );
  NOR23 U445 ( .A(n68), .B(n102), .Q(n3) );
  NAND20 U446 ( .A(n830), .B(n161), .Q(n18) );
  OAI211 U447 ( .A(n147), .B(n821), .C(n150), .Q(n146) );
  NAND20 U448 ( .A(n813), .B(n118), .Q(n13) );
  OAI211 U450 ( .A(n118), .B(n110), .C(n111), .Q(n109) );
  NAND21 U451 ( .A(A[22]), .B(B[22]), .Q(n118) );
  INV3 U452 ( .A(n199), .Q(n828) );
  NOR22 U453 ( .A(B[12]), .B(A[12]), .Q(n199) );
  NAND21 U454 ( .A(n190), .B(n832), .Q(n181) );
  INV3 U455 ( .A(n190), .Q(n829) );
  NAND21 U456 ( .A(A[20]), .B(B[20]), .Q(n132) );
  XNR22 U459 ( .A(n10), .B(n94), .Q(SUM[25]) );
  AOI211 U460 ( .A(n826), .B(n145), .C(n146), .Q(n144) );
  NOR22 U461 ( .A(n92), .B(n99), .Q(n86) );
  NOR21 U462 ( .A(B[24]), .B(A[24]), .Q(n99) );
  INV1 U463 ( .A(n160), .Q(n830) );
  NAND22 U464 ( .A(n825), .B(n145), .Q(n143) );
  NOR21 U465 ( .A(n147), .B(n823), .Q(n145) );
  NAND24 U467 ( .A(n483), .B(n484), .Q(SUM[21]) );
  XNR22 U468 ( .A(n13), .B(n119), .Q(SUM[22]) );
  OAI211 U469 ( .A(n150), .B(n140), .C(n141), .Q(n139) );
  NOR23 U470 ( .A(n140), .B(n147), .Q(n138) );
  INV0 U471 ( .A(n140), .Q(n818) );
  NOR22 U474 ( .A(B[19]), .B(A[19]), .Q(n140) );
  INV3 U475 ( .A(n130), .Q(n781) );
  AOI211 U476 ( .A(n809), .B(n77), .C(n78), .Q(n76) );
  CLKIN3 U477 ( .A(n87), .Q(n806) );
  NAND21 U478 ( .A(B[13]), .B(A[13]), .Q(n197) );
  NOR22 U479 ( .A(n136), .B(n170), .Q(n134) );
  NAND20 U480 ( .A(n825), .B(n154), .Q(n152) );
  CLKIN1 U481 ( .A(n2), .Q(n801) );
  NAND22 U482 ( .A(A[7]), .B(B[7]), .Q(n235) );
  NAND21 U483 ( .A(A[16]), .B(B[16]), .Q(n168) );
  NAND20 U484 ( .A(n824), .B(n179), .Q(n20) );
  NAND22 U485 ( .A(n217), .B(n205), .Q(n203) );
  INV0 U486 ( .A(n185), .Q(n832) );
  NAND22 U487 ( .A(n790), .B(n238), .Q(n29) );
  INV2 U489 ( .A(n237), .Q(n790) );
  INV2 U490 ( .A(n117), .Q(n813) );
  NAND20 U491 ( .A(A[23]), .B(B[23]), .Q(n111) );
  NOR20 U492 ( .A(B[31]), .B(A[31]), .Q(n36) );
  NAND20 U493 ( .A(A[4]), .B(B[4]), .Q(n251) );
  NAND20 U494 ( .A(A[5]), .B(B[5]), .Q(n246) );
  INV3 U495 ( .A(n103), .Q(n809) );
  AOI210 U496 ( .A(n2), .B(n52), .C(n55), .Q(n51) );
  NAND20 U497 ( .A(n841), .B(n215), .Q(n25) );
  NOR22 U498 ( .A(n178), .B(n185), .Q(n176) );
  INV0 U499 ( .A(n207), .Q(n833) );
  INV0 U500 ( .A(n131), .Q(n815) );
  NOR20 U501 ( .A(n237), .B(n234), .Q(n232) );
  OAI211 U502 ( .A(n238), .B(n234), .C(n235), .Q(n233) );
  NAND20 U503 ( .A(n812), .B(n111), .Q(n12) );
  NAND20 U504 ( .A(n808), .B(n100), .Q(n11) );
  INV0 U505 ( .A(n178), .Q(n824) );
  INV0 U506 ( .A(n147), .Q(n819) );
  NAND20 U507 ( .A(n819), .B(n150), .Q(n17) );
  NAND20 U508 ( .A(n840), .B(n129), .Q(n14) );
  NAND20 U509 ( .A(n52), .B(n795), .Q(n43) );
  NAND20 U510 ( .A(A[19]), .B(B[19]), .Q(n141) );
  NOR20 U511 ( .A(B[6]), .B(A[6]), .Q(n237) );
  NAND20 U512 ( .A(A[27]), .B(B[27]), .Q(n73) );
  NOR21 U513 ( .A(B[26]), .B(A[26]), .Q(n79) );
  NOR20 U514 ( .A(B[28]), .B(A[28]), .Q(n63) );
  NAND20 U515 ( .A(A[28]), .B(B[28]), .Q(n64) );
  NOR21 U516 ( .A(B[27]), .B(A[27]), .Q(n72) );
  NAND20 U517 ( .A(A[30]), .B(B[30]), .Q(n48) );
  NAND20 U518 ( .A(A[25]), .B(B[25]), .Q(n93) );
  NAND20 U519 ( .A(A[29]), .B(B[29]), .Q(n57) );
  NOR20 U520 ( .A(B[30]), .B(A[30]), .Q(n47) );
  INV3 U521 ( .A(n170), .Q(n825) );
  INV3 U522 ( .A(n8), .Q(n799) );
  NAND22 U523 ( .A(n14), .B(n130), .Q(n483) );
  NAND22 U524 ( .A(n839), .B(n781), .Q(n484) );
  INV3 U525 ( .A(n14), .Q(n839) );
  NAND22 U526 ( .A(n154), .B(n138), .Q(n136) );
  NAND22 U527 ( .A(n3), .B(n798), .Q(n59) );
  NAND20 U528 ( .A(n3), .B(n794), .Q(n39) );
  NAND22 U529 ( .A(n810), .B(n808), .Q(n95) );
  INV0 U530 ( .A(n123), .Q(n817) );
  INV3 U531 ( .A(n403), .Q(n838) );
  NAND22 U532 ( .A(n841), .B(n217), .Q(n403) );
  INV3 U533 ( .A(n240), .Q(n778) );
  INV3 U534 ( .A(n262), .Q(n776) );
  INV3 U535 ( .A(n253), .Q(n777) );
  NAND22 U536 ( .A(n833), .B(n208), .Q(n24) );
  XOR21 U537 ( .A(n26), .B(n225), .Q(SUM[9]) );
  INV0 U538 ( .A(n223), .Q(n842) );
  NAND22 U539 ( .A(n828), .B(n200), .Q(n23) );
  NAND22 U540 ( .A(n798), .B(n64), .Q(n7) );
  INV3 U541 ( .A(n3), .Q(n802) );
  NAND22 U542 ( .A(n796), .B(n57), .Q(n6) );
  INV3 U543 ( .A(n56), .Q(n796) );
  NAND22 U544 ( .A(n795), .B(n48), .Q(n5) );
  INV3 U545 ( .A(n122), .Q(n816) );
  NAND22 U546 ( .A(n803), .B(n82), .Q(n9) );
  XOR21 U547 ( .A(n778), .B(n29), .Q(SUM[6]) );
  NAND22 U548 ( .A(n804), .B(n93), .Q(n10) );
  INV3 U549 ( .A(n92), .Q(n804) );
  XNR21 U550 ( .A(n28), .B(n236), .Q(SUM[7]) );
  NAND22 U551 ( .A(n834), .B(n235), .Q(n28) );
  INV2 U552 ( .A(n234), .Q(n834) );
  NAND22 U553 ( .A(n815), .B(n132), .Q(n15) );
  NAND20 U554 ( .A(n122), .B(n813), .Q(n113) );
  XNR21 U555 ( .A(n18), .B(n162), .Q(SUM[17]) );
  XNR21 U556 ( .A(n19), .B(n169), .Q(SUM[16]) );
  AOI211 U557 ( .A(n2), .B(n798), .C(n797), .Q(n60) );
  INV3 U558 ( .A(n64), .Q(n797) );
  AOI210 U559 ( .A(n2), .B(n794), .C(n792), .Q(n40) );
  INV3 U560 ( .A(n44), .Q(n792) );
  AOI211 U561 ( .A(n55), .B(n795), .C(n793), .Q(n44) );
  INV3 U562 ( .A(n48), .Q(n793) );
  AOI210 U563 ( .A(n123), .B(n813), .C(n814), .Q(n114) );
  INV3 U564 ( .A(n118), .Q(n814) );
  NAND22 U565 ( .A(n800), .B(n73), .Q(n8) );
  INV3 U566 ( .A(n72), .Q(n800) );
  AOI210 U567 ( .A(n191), .B(n832), .C(n831), .Q(n182) );
  AOI211 U568 ( .A(n809), .B(n808), .C(n807), .Q(n96) );
  INV3 U569 ( .A(n128), .Q(n840) );
  NAND22 U570 ( .A(n812), .B(n813), .Q(n404) );
  INV3 U571 ( .A(n63), .Q(n798) );
  INV3 U572 ( .A(n99), .Q(n808) );
  INV3 U573 ( .A(n110), .Q(n812) );
  INV3 U574 ( .A(n228), .Q(n837) );
  INV3 U575 ( .A(n229), .Q(n835) );
  INV3 U576 ( .A(n43), .Q(n794) );
  XOR21 U577 ( .A(n30), .B(n247), .Q(SUM[5]) );
  NAND22 U578 ( .A(n789), .B(n246), .Q(n30) );
  AOI211 U579 ( .A(n777), .B(n787), .C(n786), .Q(n247) );
  XOR21 U580 ( .A(n33), .B(n776), .Q(SUM[2]) );
  NAND22 U581 ( .A(n784), .B(n260), .Q(n33) );
  INV3 U582 ( .A(n259), .Q(n784) );
  XOR21 U583 ( .A(n266), .B(n34), .Q(SUM[1]) );
  NAND22 U584 ( .A(n783), .B(n264), .Q(n34) );
  INV3 U585 ( .A(n263), .Q(n783) );
  NAND22 U586 ( .A(n787), .B(n789), .Q(n241) );
  AOI211 U587 ( .A(n789), .B(n786), .C(n788), .Q(n242) );
  INV3 U588 ( .A(n246), .Q(n788) );
  XNR21 U589 ( .A(n32), .B(n258), .Q(SUM[3]) );
  NAND22 U590 ( .A(n785), .B(n257), .Q(n32) );
  INV3 U591 ( .A(n256), .Q(n785) );
  AOI211 U592 ( .A(n262), .B(n254), .C(n255), .Q(n253) );
  NOR21 U593 ( .A(n256), .B(n259), .Q(n254) );
  XNR21 U594 ( .A(n31), .B(n777), .Q(SUM[4]) );
  NAND22 U595 ( .A(n787), .B(n251), .Q(n31) );
  INV3 U596 ( .A(n251), .Q(n786) );
  XNR21 U597 ( .A(n4), .B(n38), .Q(SUM[31]) );
  NAND22 U598 ( .A(n791), .B(n37), .Q(n4) );
  NAND22 U599 ( .A(A[31]), .B(B[31]), .Q(n37) );
  NOR22 U600 ( .A(B[18]), .B(A[18]), .Q(n147) );
  NOR22 U601 ( .A(B[15]), .B(A[15]), .Q(n178) );
  NOR21 U602 ( .A(B[20]), .B(A[20]), .Q(n131) );
  NAND21 U603 ( .A(A[18]), .B(B[18]), .Q(n150) );
  NAND21 U604 ( .A(A[21]), .B(B[21]), .Q(n129) );
  INV3 U605 ( .A(n47), .Q(n795) );
  INV3 U606 ( .A(n36), .Q(n791) );
  NAND20 U607 ( .A(A[6]), .B(B[6]), .Q(n238) );
  INV3 U608 ( .A(n245), .Q(n789) );
  NOR20 U609 ( .A(B[5]), .B(A[5]), .Q(n245) );
  INV3 U610 ( .A(n35), .Q(SUM[0]) );
  NAND22 U611 ( .A(n775), .B(n266), .Q(n35) );
  INV3 U612 ( .A(n265), .Q(n775) );
  NOR20 U613 ( .A(B[0]), .B(A[0]), .Q(n265) );
  INV3 U614 ( .A(n250), .Q(n787) );
  NOR20 U615 ( .A(B[4]), .B(A[4]), .Q(n250) );
  NOR20 U616 ( .A(B[3]), .B(A[3]), .Q(n256) );
  NOR20 U617 ( .A(B[2]), .B(A[2]), .Q(n259) );
  NAND20 U618 ( .A(A[0]), .B(B[0]), .Q(n266) );
  NAND20 U619 ( .A(A[2]), .B(B[2]), .Q(n260) );
  NOR20 U620 ( .A(B[1]), .B(A[1]), .Q(n263) );
  NAND20 U621 ( .A(A[1]), .B(B[1]), .Q(n264) );
  NAND20 U622 ( .A(A[3]), .B(B[3]), .Q(n257) );
  INV2 U623 ( .A(n191), .Q(n827) );
endmodule


module adder_28 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_28_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_27_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n265, n266, n268, n269, n270, n271, n272, n273,
         n274, n275, n277, n278, n279, n280, n281, n416, n427, n582, n584,
         n585, n589, n660, n662, n735, n741, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n880, n881, n882;

  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U207 ( .A(n188), .B(n871), .C(n189), .Q(n187) );
  OAI212 U219 ( .A(n197), .B(n871), .C(n198), .Q(n196) );
  OAI212 U227 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  OAI212 U233 ( .A(n208), .B(n871), .C(n209), .Q(n207) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n223), .B(n231), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n871), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n868), .B(n871), .C(n866), .Q(n232) );
  OAI212 U281 ( .A(n244), .B(n871), .C(n245), .Q(n243) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U298 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n881), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U465 ( .A(n817), .B(n82), .C(n83), .Q(n81) );
  OAI212 U494 ( .A(n152), .B(n113), .C(n114), .Q(n112) );
  OAI212 U484 ( .A(n817), .B(n120), .C(n121), .Q(n119) );
  OAI212 U416 ( .A(n73), .B(n817), .C(n74), .Q(n72) );
  OAI212 U458 ( .A(n851), .B(n817), .C(n849), .Q(n164) );
  OAI212 U438 ( .A(n158), .B(n817), .C(n159), .Q(n157) );
  OAI212 U426 ( .A(n42), .B(n817), .C(n43), .Q(n41) );
  OAI212 U429 ( .A(n91), .B(n817), .C(n92), .Q(n90) );
  OAI212 U452 ( .A(n177), .B(n173), .C(n808), .Q(n662) );
  OAI212 U459 ( .A(n176), .B(n817), .C(n177), .Q(n175) );
  OAI212 U487 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U499 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  AOI212 U509 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U434 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U440 ( .A(n151), .B(n817), .C(n660), .Q(n146) );
  OAI212 U444 ( .A(n837), .B(n817), .C(n835), .Q(n108) );
  OAI212 U445 ( .A(n102), .B(n817), .C(n103), .Q(n101) );
  OAI212 U449 ( .A(n129), .B(n817), .C(n130), .Q(n128) );
  OAI212 U512 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U528 ( .A(n256), .B(n416), .C(n253), .Q(n251) );
  CLKIN3 U349 ( .A(n151), .Q(n846) );
  NAND21 U350 ( .A(n111), .B(n66), .Q(n64) );
  NAND23 U351 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NAND21 U352 ( .A(A[17]), .B(B[17]), .Q(n808) );
  NAND20 U353 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NAND24 U354 ( .A(n153), .B(n171), .Q(n151) );
  NOR23 U355 ( .A(n144), .B(n137), .Q(n135) );
  NOR23 U356 ( .A(n809), .B(A[21]), .Q(n137) );
  CLKIN1 U357 ( .A(n832), .Q(n810) );
  INV2 U358 ( .A(n98), .Q(n832) );
  NOR24 U359 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR24 U360 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR23 U361 ( .A(B[12]), .B(A[12]), .Q(n212) );
  INV2 U362 ( .A(n46), .Q(n819) );
  NOR24 U363 ( .A(A[25]), .B(B[25]), .Q(n99) );
  NAND23 U364 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND24 U365 ( .A(n111), .B(n828), .Q(n584) );
  NAND26 U366 ( .A(n135), .B(n741), .Q(n113) );
  NOR24 U367 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR24 U368 ( .A(n185), .B(n194), .Q(n183) );
  NOR24 U369 ( .A(B[15]), .B(A[15]), .Q(n185) );
  INV1 U370 ( .A(n220), .Q(n858) );
  NOR22 U371 ( .A(n162), .B(n155), .Q(n153) );
  NOR22 U372 ( .A(n117), .B(n126), .Q(n741) );
  NOR22 U373 ( .A(A[18]), .B(B[18]), .Q(n162) );
  NOR23 U374 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR23 U375 ( .A(n824), .B(n584), .Q(n585) );
  NOR22 U376 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR22 U377 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NOR23 U378 ( .A(B[13]), .B(A[13]), .Q(n205) );
  BUF2 U379 ( .A(n127), .Q(n816) );
  NAND22 U380 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND22 U381 ( .A(A[24]), .B(B[24]), .Q(n107) );
  XOR21 U382 ( .A(n22), .B(n817), .Q(SUM[16]) );
  INV3 U383 ( .A(n163), .Q(n847) );
  BUF6 U384 ( .A(B[21]), .Q(n809) );
  NAND22 U385 ( .A(n80), .B(n827), .Q(n11) );
  OAI211 U386 ( .A(n88), .B(n832), .C(n89), .Q(n85) );
  CLKIN1 U387 ( .A(n839), .Q(n814) );
  INV3 U388 ( .A(n88), .Q(n829) );
  INV2 U389 ( .A(n826), .Q(n811) );
  INV3 U390 ( .A(n811), .Q(n812) );
  BUF15 U391 ( .A(n112), .Q(n813) );
  XNR22 U392 ( .A(n19), .B(n157), .Q(SUM[19]) );
  XNR22 U393 ( .A(n18), .B(n146), .Q(SUM[20]) );
  CLKIN3 U394 ( .A(n117), .Q(n836) );
  XNR22 U395 ( .A(n20), .B(n164), .Q(SUM[18]) );
  AOI211 U396 ( .A(n844), .B(n135), .C(n814), .Q(n130) );
  NOR23 U397 ( .A(n46), .B(n6), .Q(n44) );
  INV0 U398 ( .A(n185), .Q(n853) );
  NAND23 U399 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NOR23 U400 ( .A(n205), .B(n212), .Q(n203) );
  XNR22 U401 ( .A(n21), .B(n175), .Q(SUM[17]) );
  INV2 U402 ( .A(n135), .Q(n841) );
  NAND28 U403 ( .A(n735), .B(n156), .Q(n154) );
  NAND22 U404 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND23 U405 ( .A(n427), .B(n822), .Q(n56) );
  AOI212 U406 ( .A(n813), .B(n828), .C(n812), .Q(n74) );
  NOR23 U407 ( .A(n99), .B(n106), .Q(n97) );
  NOR23 U408 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND21 U409 ( .A(A[21]), .B(n809), .Q(n138) );
  NOR23 U410 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR22 U411 ( .A(n70), .B(n6), .Q(n66) );
  CLKIN6 U412 ( .A(n6), .Q(n828) );
  XNR22 U413 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND21 U414 ( .A(A[25]), .B(B[25]), .Q(n100) );
  INV2 U415 ( .A(n813), .Q(n835) );
  OAI212 U417 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  NAND28 U418 ( .A(n97), .B(n77), .Q(n6) );
  NAND21 U419 ( .A(A[29]), .B(B[29]), .Q(n62) );
  XNR22 U420 ( .A(n15), .B(n119), .Q(SUM[23]) );
  AOI212 U421 ( .A(n813), .B(n66), .C(n67), .Q(n65) );
  AOI212 U422 ( .A(n98), .B(n77), .C(n78), .Q(n815) );
  NAND22 U423 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NOR24 U424 ( .A(A[22]), .B(B[22]), .Q(n126) );
  NOR21 U425 ( .A(n824), .B(n6), .Q(n55) );
  NAND24 U427 ( .A(n585), .B(n854), .Q(n589) );
  INV10 U428 ( .A(n817), .Q(n854) );
  BUF15 U430 ( .A(n178), .Q(n817) );
  NAND22 U431 ( .A(n826), .B(n59), .Q(n427) );
  INV2 U432 ( .A(n136), .Q(n839) );
  OAI212 U433 ( .A(n140), .B(n817), .C(n141), .Q(n139) );
  XNR22 U435 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U436 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND21 U437 ( .A(B[23]), .B(A[23]), .Q(n118) );
  NAND21 U439 ( .A(n100), .B(n830), .Q(n13) );
  NAND23 U441 ( .A(n582), .B(n47), .Q(n45) );
  AOI212 U442 ( .A(n153), .B(n662), .C(n154), .Q(n660) );
  XNR22 U443 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U446 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NAND21 U447 ( .A(n846), .B(n135), .Q(n129) );
  OAI210 U448 ( .A(n194), .B(n861), .C(n195), .Q(n191) );
  AOI211 U450 ( .A(n844), .B(n843), .C(n842), .Q(n141) );
  INV3 U451 ( .A(n144), .Q(n843) );
  AOI212 U453 ( .A(n813), .B(n97), .C(n810), .Q(n92) );
  XNR22 U454 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND24 U455 ( .A(n589), .B(n54), .Q(n52) );
  AOI212 U456 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND21 U457 ( .A(n111), .B(n828), .Q(n73) );
  NAND21 U460 ( .A(n111), .B(n84), .Q(n82) );
  NAND21 U461 ( .A(n111), .B(n44), .Q(n42) );
  NAND21 U462 ( .A(n111), .B(n833), .Q(n102) );
  NAND21 U463 ( .A(n111), .B(n97), .Q(n91) );
  INV2 U464 ( .A(n111), .Q(n837) );
  OAI211 U466 ( .A(n126), .B(n839), .C(n816), .Q(n123) );
  OAI210 U467 ( .A(n219), .B(n871), .C(n220), .Q(n214) );
  CLKIN6 U468 ( .A(n5), .Q(n826) );
  XNR22 U469 ( .A(n9), .B(n63), .Q(SUM[29]) );
  OAI212 U470 ( .A(n817), .B(n64), .C(n65), .Q(n63) );
  INV0 U471 ( .A(n107), .Q(n834) );
  XNR22 U472 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U473 ( .A(n17), .B(n139), .Q(SUM[21]) );
  AOI212 U474 ( .A(n813), .B(n84), .C(n85), .Q(n83) );
  AOI212 U475 ( .A(n813), .B(n833), .C(n834), .Q(n103) );
  AOI212 U476 ( .A(n813), .B(n55), .C(n56), .Q(n54) );
  NOR24 U477 ( .A(n61), .B(n70), .Q(n59) );
  INV2 U478 ( .A(n70), .Q(n825) );
  NOR24 U479 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR21 U480 ( .A(n126), .B(n841), .Q(n122) );
  OAI212 U481 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  NAND21 U482 ( .A(B[27]), .B(A[27]), .Q(n80) );
  NOR24 U483 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND22 U485 ( .A(A[15]), .B(B[15]), .Q(n186) );
  INV0 U486 ( .A(n79), .Q(n827) );
  INV2 U488 ( .A(n126), .Q(n838) );
  NOR22 U489 ( .A(n117), .B(n126), .Q(n115) );
  NOR24 U490 ( .A(n113), .B(n151), .Q(n111) );
  NOR24 U491 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR24 U492 ( .A(n79), .B(n88), .Q(n77) );
  NAND20 U493 ( .A(n833), .B(n107), .Q(n14) );
  INV2 U495 ( .A(n106), .Q(n833) );
  NAND24 U496 ( .A(n203), .B(n183), .Q(n181) );
  XNR22 U497 ( .A(n10), .B(n72), .Q(SUM[28]) );
  INV1 U498 ( .A(n162), .Q(n848) );
  NOR23 U500 ( .A(n173), .B(n176), .Q(n171) );
  NAND22 U501 ( .A(n171), .B(n848), .Q(n158) );
  INV1 U502 ( .A(n171), .Q(n851) );
  INV0 U503 ( .A(n137), .Q(n840) );
  NAND22 U504 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U505 ( .A(n864), .B(n213), .Q(n26) );
  CLKIN3 U506 ( .A(n204), .Q(n861) );
  INV0 U507 ( .A(n99), .Q(n830) );
  AOI212 U508 ( .A(n813), .B(n44), .C(n45), .Q(n43) );
  INV2 U510 ( .A(n97), .Q(n831) );
  INV3 U511 ( .A(n59), .Q(n824) );
  NAND23 U513 ( .A(n59), .B(n820), .Q(n46) );
  NAND21 U514 ( .A(n845), .B(n156), .Q(n19) );
  NAND20 U515 ( .A(n848), .B(n163), .Q(n20) );
  NAND22 U516 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NOR23 U517 ( .A(n88), .B(n831), .Q(n84) );
  NOR24 U518 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND24 U519 ( .A(n847), .B(n845), .Q(n735) );
  AOI212 U520 ( .A(n115), .B(n136), .C(n116), .Q(n114) );
  OAI212 U521 ( .A(n137), .B(n145), .C(n138), .Q(n136) );
  AOI212 U522 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  NAND23 U523 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND22 U524 ( .A(A[18]), .B(B[18]), .Q(n163) );
  AOI211 U525 ( .A(n844), .B(n122), .C(n123), .Q(n121) );
  NAND21 U526 ( .A(n846), .B(n122), .Q(n120) );
  NAND21 U527 ( .A(n846), .B(n843), .Q(n140) );
  CLKIN1 U529 ( .A(n60), .Q(n822) );
  INV0 U530 ( .A(n145), .Q(n842) );
  NAND21 U531 ( .A(n869), .B(n245), .Q(n30) );
  NAND20 U532 ( .A(n857), .B(n203), .Q(n197) );
  AOI211 U533 ( .A(n60), .B(n820), .C(n821), .Q(n47) );
  INV2 U534 ( .A(n51), .Q(n821) );
  INV0 U535 ( .A(n212), .Q(n864) );
  CLKIN0 U536 ( .A(n231), .Q(n859) );
  INV2 U537 ( .A(n230), .Q(n860) );
  INV2 U538 ( .A(n244), .Q(n869) );
  NOR20 U539 ( .A(n241), .B(n244), .Q(n239) );
  NOR20 U540 ( .A(n416), .B(n255), .Q(n250) );
  NAND21 U541 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND20 U542 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND20 U543 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR22 U544 ( .A(n181), .B(n219), .Q(n179) );
  AOI210 U545 ( .A(n858), .B(n203), .C(n204), .Q(n198) );
  NAND20 U546 ( .A(n857), .B(n190), .Q(n188) );
  AOI211 U547 ( .A(n858), .B(n190), .C(n191), .Q(n189) );
  NAND20 U548 ( .A(n860), .B(n231), .Q(n28) );
  NAND20 U549 ( .A(n224), .B(n856), .Q(n27) );
  NOR20 U550 ( .A(A[10]), .B(B[10]), .Q(n230) );
  NAND20 U551 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND21 U552 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U553 ( .A(n39), .Q(n818) );
  NAND21 U554 ( .A(n62), .B(n823), .Q(n9) );
  INV3 U555 ( .A(n660), .Q(n844) );
  INV3 U556 ( .A(n219), .Q(n857) );
  INV0 U557 ( .A(n662), .Q(n849) );
  AOI210 U558 ( .A(n662), .B(n848), .C(n847), .Q(n159) );
  INV3 U559 ( .A(n203), .Q(n863) );
  AOI211 U560 ( .A(n877), .B(n258), .C(n259), .Q(n257) );
  NAND22 U561 ( .A(n239), .B(n221), .Q(n219) );
  INV3 U562 ( .A(n247), .Q(n871) );
  INV3 U563 ( .A(n268), .Q(n877) );
  NAND22 U564 ( .A(n239), .B(n860), .Q(n226) );
  INV3 U565 ( .A(n240), .Q(n866) );
  INV3 U566 ( .A(n239), .Q(n868) );
  NOR21 U567 ( .A(n194), .B(n863), .Q(n190) );
  NAND22 U568 ( .A(n857), .B(n864), .Q(n208) );
  AOI210 U569 ( .A(n858), .B(n864), .C(n865), .Q(n209) );
  INV3 U570 ( .A(n213), .Q(n865) );
  AOI211 U571 ( .A(n240), .B(n860), .C(n859), .Q(n227) );
  INV3 U572 ( .A(n155), .Q(n845) );
  NAND22 U573 ( .A(n826), .B(n819), .Q(n582) );
  INV3 U574 ( .A(n223), .Q(n856) );
  INV3 U575 ( .A(n61), .Q(n823) );
  INV3 U576 ( .A(n173), .Q(n850) );
  INV3 U577 ( .A(n265), .Q(n873) );
  INV3 U578 ( .A(n194), .Q(n855) );
  INV3 U579 ( .A(n176), .Q(n852) );
  INV3 U580 ( .A(n205), .Q(n862) );
  NAND22 U581 ( .A(n867), .B(n242), .Q(n29) );
  INV3 U582 ( .A(n241), .Q(n867) );
  NAND22 U583 ( .A(n872), .B(n253), .Q(n31) );
  INV3 U584 ( .A(n416), .Q(n872) );
  NAND22 U585 ( .A(n875), .B(n261), .Q(n33) );
  INV3 U586 ( .A(n260), .Q(n875) );
  INV3 U587 ( .A(n255), .Q(n870) );
  INV3 U588 ( .A(n278), .Q(n882) );
  NAND22 U589 ( .A(n878), .B(n272), .Q(n35) );
  INV3 U590 ( .A(n271), .Q(n878) );
  INV3 U591 ( .A(n274), .Q(n876) );
  AOI211 U592 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U593 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U594 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U595 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U596 ( .A(n223), .B(n230), .Q(n221) );
  NOR21 U597 ( .A(n260), .B(n265), .Q(n258) );
  INV3 U598 ( .A(n277), .Q(n881) );
  INV3 U599 ( .A(n266), .Q(n874) );
  NOR21 U600 ( .A(B[7]), .B(A[7]), .Q(n416) );
  NOR21 U601 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NOR21 U602 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR21 U603 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR21 U604 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U605 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U606 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U607 ( .A(B[11]), .B(A[11]), .Q(n224) );
  INV3 U608 ( .A(n50), .Q(n820) );
  NOR21 U609 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NOR21 U610 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U611 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND22 U612 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U613 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U614 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND22 U615 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U616 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND22 U617 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND22 U618 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NOR21 U619 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U620 ( .A(n280), .Q(n880) );
  NOR21 U621 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U622 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U623 ( .A(n816), .B(n838), .Q(n16) );
  NAND22 U624 ( .A(n818), .B(n40), .Q(n7) );
  NAND20 U625 ( .A(n808), .B(n850), .Q(n21) );
  NAND20 U626 ( .A(n843), .B(n145), .Q(n18) );
  NAND20 U627 ( .A(n836), .B(n118), .Q(n15) );
  NAND20 U628 ( .A(n829), .B(n89), .Q(n12) );
  NAND20 U629 ( .A(n825), .B(n71), .Q(n10) );
  NAND20 U630 ( .A(n852), .B(n177), .Q(n22) );
  XNR21 U631 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U632 ( .A(n195), .B(n855), .Q(n24) );
  XNR21 U633 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U634 ( .A(n862), .B(n206), .Q(n25) );
  XNR21 U635 ( .A(n27), .B(n225), .Q(SUM[11]) );
  XOR21 U636 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U637 ( .A(n877), .B(n873), .C(n874), .Q(n262) );
  XOR21 U638 ( .A(n30), .B(n871), .Q(SUM[8]) );
  NAND20 U639 ( .A(n820), .B(n51), .Q(n8) );
  NAND20 U640 ( .A(n840), .B(n138), .Q(n17) );
  XNR21 U641 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U642 ( .A(n853), .B(n186), .Q(n23) );
  XNR21 U643 ( .A(n26), .B(n214), .Q(SUM[12]) );
  XOR21 U644 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND22 U645 ( .A(n870), .B(n256), .Q(n32) );
  XNR21 U646 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XNR21 U647 ( .A(n34), .B(n877), .Q(SUM[4]) );
  NAND22 U648 ( .A(n873), .B(n266), .Q(n34) );
  XNR21 U649 ( .A(n29), .B(n243), .Q(SUM[9]) );
  XNR21 U650 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XOR21 U651 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U652 ( .A(n882), .B(n279), .Q(n37) );
  XOR21 U653 ( .A(n36), .B(n881), .Q(SUM[2]) );
  NAND22 U654 ( .A(n876), .B(n275), .Q(n36) );
  XNR21 U655 ( .A(n35), .B(n273), .Q(SUM[3]) );
  INV3 U656 ( .A(n38), .Q(SUM[0]) );
  NAND22 U657 ( .A(n880), .B(n281), .Q(n38) );
  OAI211 U658 ( .A(n815), .B(n70), .C(n71), .Q(n67) );
endmodule


module adder_27 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_27_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_26_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n420, n421,
         n430, n436, n437, n658, n665, n666, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U306 ( .A(n260), .B(n266), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  AOI212 U488 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U489 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  AOI212 U507 ( .A(n247), .B(n179), .C(n810), .Q(n178) );
  OAI212 U467 ( .A(n102), .B(n831), .C(n103), .Q(n101) );
  OAI212 U472 ( .A(n91), .B(n831), .C(n92), .Q(n90) );
  OAI212 U473 ( .A(n82), .B(n831), .C(n83), .Q(n81) );
  OAI212 U665 ( .A(n248), .B(n268), .C(n249), .Q(n420) );
  OAI212 U411 ( .A(n163), .B(n809), .C(n156), .Q(n154) );
  OAI212 U431 ( .A(n127), .B(n832), .C(n118), .Q(n116) );
  OAI212 U447 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U455 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U466 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  OAI212 U470 ( .A(n241), .B(n245), .C(n242), .Q(n240) );
  OAI212 U509 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U656 ( .A(n185), .B(n195), .C(n186), .Q(n184) );
  OAI212 U521 ( .A(n64), .B(n831), .C(n65), .Q(n63) );
  OAI212 U659 ( .A(n274), .B(n884), .C(n275), .Q(n273) );
  OAI212 U391 ( .A(n53), .B(n831), .C(n54), .Q(n52) );
  OAI212 U460 ( .A(n73), .B(n831), .C(n74), .Q(n72) );
  OAI212 U420 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U422 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI212 U423 ( .A(n837), .B(n5), .C(n838), .Q(n56) );
  OAI212 U443 ( .A(n248), .B(n811), .C(n249), .Q(n247) );
  OAI212 U501 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U349 ( .A(n158), .B(n813), .C(n159), .Q(n157) );
  INV2 U350 ( .A(n152), .Q(n857) );
  INV6 U351 ( .A(n101), .Q(n817) );
  INV0 U352 ( .A(n871), .Q(n807) );
  INV4 U353 ( .A(n220), .Q(n871) );
  NOR22 U354 ( .A(n260), .B(n265), .Q(n258) );
  AOI211 U355 ( .A(n871), .B(n190), .C(n191), .Q(n189) );
  OAI212 U356 ( .A(n176), .B(n178), .C(n177), .Q(n175) );
  NAND22 U357 ( .A(n111), .B(n66), .Q(n64) );
  NOR21 U358 ( .A(n181), .B(n219), .Q(n658) );
  NAND28 U359 ( .A(n203), .B(n183), .Q(n181) );
  XNR22 U360 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XNR22 U361 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NOR22 U362 ( .A(n173), .B(n176), .Q(n171) );
  INV3 U363 ( .A(n155), .Q(n808) );
  INV6 U364 ( .A(n808), .Q(n809) );
  CLKIN2 U365 ( .A(n128), .Q(n821) );
  OAI211 U366 ( .A(n129), .B(n178), .C(n130), .Q(n128) );
  XNR22 U367 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NOR23 U368 ( .A(n79), .B(n88), .Q(n77) );
  XNR22 U369 ( .A(n23), .B(n187), .Q(SUM[15]) );
  XNR22 U370 ( .A(n225), .B(n27), .Q(SUM[11]) );
  NAND20 U371 ( .A(n171), .B(n858), .Q(n158) );
  INV0 U372 ( .A(n171), .Q(n864) );
  NAND24 U373 ( .A(n171), .B(n153), .Q(n151) );
  INV3 U374 ( .A(n97), .Q(n845) );
  NAND21 U375 ( .A(n111), .B(n97), .Q(n91) );
  AOI212 U376 ( .A(n815), .B(n97), .C(n98), .Q(n92) );
  NAND23 U377 ( .A(n97), .B(n77), .Q(n6) );
  NOR23 U378 ( .A(n99), .B(n106), .Q(n97) );
  NAND24 U379 ( .A(n135), .B(n115), .Q(n113) );
  CLKIN6 U380 ( .A(n135), .Q(n855) );
  NAND20 U381 ( .A(n859), .B(n135), .Q(n129) );
  NOR23 U382 ( .A(n137), .B(n144), .Q(n135) );
  AOI211 U383 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  BUF12 U384 ( .A(n421), .Q(n831) );
  AOI211 U385 ( .A(n420), .B(n658), .C(n437), .Q(n421) );
  NOR22 U386 ( .A(n252), .B(n255), .Q(n250) );
  NOR21 U387 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U388 ( .A(n258), .B(n250), .Q(n248) );
  NOR22 U389 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR21 U390 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR21 U392 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND22 U393 ( .A(n871), .B(n868), .Q(n436) );
  NOR21 U394 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR22 U395 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR21 U396 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR21 U397 ( .A(n837), .B(n6), .Q(n55) );
  NAND22 U398 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR21 U399 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR22 U400 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND23 U401 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR23 U402 ( .A(A[13]), .B(B[13]), .Q(n205) );
  NAND22 U403 ( .A(n870), .B(n896), .Q(n208) );
  NOR23 U404 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR21 U405 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NAND22 U406 ( .A(n826), .B(n827), .Q(SUM[21]) );
  NAND22 U407 ( .A(n825), .B(n824), .Q(n827) );
  BUF12 U408 ( .A(n180), .Q(n810) );
  OAI211 U409 ( .A(n140), .B(n178), .C(n141), .Q(n139) );
  INV3 U410 ( .A(n829), .Q(n886) );
  AOI212 U412 ( .A(n277), .B(n269), .C(n270), .Q(n811) );
  NOR24 U413 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NOR22 U414 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NAND21 U415 ( .A(n854), .B(n145), .Q(n18) );
  NAND21 U416 ( .A(A[3]), .B(B[3]), .Q(n272) );
  AOI212 U417 ( .A(n247), .B(n179), .C(n810), .Q(n812) );
  AOI212 U418 ( .A(n247), .B(n179), .C(n810), .Q(n813) );
  CLKIN0 U419 ( .A(n213), .Q(n897) );
  NOR24 U421 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NAND22 U424 ( .A(n111), .B(n848), .Q(n102) );
  NOR23 U425 ( .A(n113), .B(n151), .Q(n111) );
  NOR22 U426 ( .A(B[23]), .B(A[23]), .Q(n117) );
  CLKIN6 U427 ( .A(n112), .Q(n814) );
  INV8 U428 ( .A(n814), .Q(n815) );
  OAI210 U429 ( .A(n42), .B(n831), .C(n43), .Q(n41) );
  INV2 U430 ( .A(n139), .Q(n825) );
  NOR23 U432 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND22 U433 ( .A(B[5]), .B(A[5]), .Q(n261) );
  INV0 U434 ( .A(n173), .Q(n863) );
  INV3 U435 ( .A(n162), .Q(n858) );
  NOR21 U436 ( .A(n194), .B(n894), .Q(n190) );
  AOI211 U437 ( .A(n857), .B(n135), .C(n136), .Q(n130) );
  AOI211 U438 ( .A(n815), .B(n55), .C(n56), .Q(n54) );
  AOI212 U439 ( .A(n815), .B(n848), .C(n847), .Q(n103) );
  AOI211 U440 ( .A(n815), .B(n841), .C(n842), .Q(n74) );
  AOI211 U441 ( .A(n815), .B(n66), .C(n67), .Q(n65) );
  AOI212 U442 ( .A(n815), .B(n84), .C(n85), .Q(n83) );
  NOR23 U444 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR24 U445 ( .A(A[15]), .B(B[15]), .Q(n185) );
  NAND22 U446 ( .A(n436), .B(n182), .Q(n437) );
  NAND20 U448 ( .A(n870), .B(n203), .Q(n197) );
  INV3 U449 ( .A(n203), .Q(n894) );
  NOR24 U450 ( .A(n181), .B(n219), .Q(n179) );
  INV2 U451 ( .A(n181), .Q(n868) );
  NAND23 U452 ( .A(n821), .B(n820), .Q(n823) );
  NOR24 U453 ( .A(n194), .B(n185), .Q(n183) );
  NAND21 U454 ( .A(n891), .B(n261), .Q(n33) );
  NAND21 U456 ( .A(A[11]), .B(B[11]), .Q(n224) );
  AOI210 U457 ( .A(n871), .B(n896), .C(n897), .Q(n209) );
  NAND22 U458 ( .A(n59), .B(n835), .Q(n46) );
  NOR24 U459 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND20 U461 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND26 U462 ( .A(n239), .B(n221), .Q(n219) );
  NAND20 U463 ( .A(n239), .B(n869), .Q(n226) );
  INV0 U464 ( .A(n239), .Q(n875) );
  NOR22 U465 ( .A(n244), .B(n241), .Q(n239) );
  NAND22 U468 ( .A(n13), .B(n101), .Q(n818) );
  NAND26 U469 ( .A(n816), .B(n817), .Q(n819) );
  NAND28 U471 ( .A(n818), .B(n819), .Q(SUM[25]) );
  INV6 U474 ( .A(n13), .Q(n816) );
  NAND21 U475 ( .A(n100), .B(n844), .Q(n13) );
  NAND22 U476 ( .A(A[6]), .B(B[6]), .Q(n256) );
  OAI212 U477 ( .A(n245), .B(n829), .C(n242), .Q(n430) );
  OAI211 U478 ( .A(n151), .B(n812), .C(n152), .Q(n146) );
  XNR22 U479 ( .A(n20), .B(n164), .Q(SUM[18]) );
  OAI211 U480 ( .A(n864), .B(n813), .C(n862), .Q(n164) );
  NAND21 U481 ( .A(n16), .B(n128), .Q(n822) );
  NAND24 U482 ( .A(n822), .B(n823), .Q(SUM[22]) );
  INV3 U483 ( .A(n16), .Q(n820) );
  NAND21 U484 ( .A(n139), .B(n17), .Q(n826) );
  INV3 U485 ( .A(n17), .Q(n824) );
  OAI212 U486 ( .A(n208), .B(n877), .C(n209), .Q(n207) );
  OAI212 U487 ( .A(n226), .B(n877), .C(n227), .Q(n225) );
  BUF2 U490 ( .A(n223), .Q(n828) );
  AOI211 U491 ( .A(n857), .B(n122), .C(n123), .Q(n121) );
  NOR23 U492 ( .A(n205), .B(n212), .Q(n203) );
  INV1 U493 ( .A(n212), .Q(n896) );
  XNR22 U494 ( .A(n214), .B(n26), .Q(SUM[12]) );
  NAND21 U495 ( .A(A[17]), .B(B[17]), .Q(n174) );
  CLKIN6 U496 ( .A(n219), .Q(n870) );
  XNR22 U497 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND22 U498 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND21 U499 ( .A(A[7]), .B(B[7]), .Q(n253) );
  CLKIN3 U500 ( .A(n430), .Q(n873) );
  AOI212 U502 ( .A(n430), .B(n869), .C(n872), .Q(n227) );
  INV1 U503 ( .A(n230), .Q(n869) );
  INV0 U504 ( .A(n194), .Q(n867) );
  XNR22 U505 ( .A(n207), .B(n25), .Q(SUM[13]) );
  NOR23 U506 ( .A(n230), .B(n223), .Q(n221) );
  BUF2 U508 ( .A(n241), .Q(n829) );
  NAND22 U510 ( .A(A[9]), .B(B[9]), .Q(n242) );
  INV0 U511 ( .A(n176), .Q(n866) );
  NAND21 U512 ( .A(B[15]), .B(A[15]), .Q(n186) );
  NAND22 U513 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NOR24 U514 ( .A(B[11]), .B(A[11]), .Q(n223) );
  XNR22 U515 ( .A(n9), .B(n63), .Q(SUM[29]) );
  INV2 U516 ( .A(n892), .Q(n830) );
  INV1 U517 ( .A(n204), .Q(n892) );
  NAND21 U518 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND21 U519 ( .A(A[26]), .B(B[26]), .Q(n89) );
  XNR22 U520 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI212 U522 ( .A(n850), .B(n831), .C(n814), .Q(n108) );
  INV0 U523 ( .A(n185), .Q(n885) );
  XNR22 U524 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NAND20 U525 ( .A(n886), .B(n242), .Q(n29) );
  NAND20 U526 ( .A(n863), .B(n174), .Q(n21) );
  OAI211 U527 ( .A(n219), .B(n877), .C(n807), .Q(n214) );
  NAND22 U528 ( .A(B[12]), .B(A[12]), .Q(n213) );
  INV6 U529 ( .A(n420), .Q(n877) );
  INV0 U530 ( .A(n205), .Q(n893) );
  OAI212 U531 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U532 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  NAND22 U533 ( .A(n870), .B(n190), .Q(n188) );
  NAND20 U534 ( .A(n876), .B(n256), .Q(n32) );
  OAI210 U535 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NAND24 U536 ( .A(n665), .B(n666), .Q(SUM[17]) );
  NAND21 U537 ( .A(A[22]), .B(B[22]), .Q(n127) );
  OAI210 U538 ( .A(n126), .B(n853), .C(n127), .Q(n123) );
  NAND20 U539 ( .A(n851), .B(n127), .Q(n16) );
  OAI211 U540 ( .A(n194), .B(n892), .C(n195), .Q(n191) );
  OAI212 U541 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  NAND22 U542 ( .A(n848), .B(n107), .Q(n14) );
  NAND21 U543 ( .A(A[24]), .B(B[24]), .Q(n107) );
  INV3 U544 ( .A(n98), .Q(n846) );
  XNR22 U545 ( .A(n10), .B(n72), .Q(SUM[28]) );
  INV0 U546 ( .A(n137), .Q(n890) );
  OAI211 U547 ( .A(n120), .B(n813), .C(n121), .Q(n119) );
  AOI212 U548 ( .A(n250), .B(n259), .C(n251), .Q(n249) );
  OAI211 U549 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NOR21 U550 ( .A(B[29]), .B(A[29]), .Q(n61) );
  OAI210 U551 ( .A(n244), .B(n877), .C(n245), .Q(n243) );
  OAI211 U552 ( .A(n197), .B(n877), .C(n198), .Q(n196) );
  OAI211 U553 ( .A(n875), .B(n877), .C(n873), .Q(n232) );
  OAI211 U554 ( .A(n188), .B(n877), .C(n189), .Q(n187) );
  XOR21 U555 ( .A(n812), .B(n22), .Q(SUM[16]) );
  XNR22 U556 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND21 U557 ( .A(A[18]), .B(B[18]), .Q(n163) );
  INV1 U558 ( .A(n6), .Q(n841) );
  OAI210 U559 ( .A(n88), .B(n846), .C(n89), .Q(n85) );
  CLKIN1 U560 ( .A(n111), .Q(n850) );
  NAND21 U561 ( .A(n841), .B(n111), .Q(n73) );
  BUF2 U562 ( .A(n117), .Q(n832) );
  INV3 U563 ( .A(n151), .Q(n859) );
  NAND22 U564 ( .A(n111), .B(n84), .Q(n82) );
  INV2 U565 ( .A(n5), .Q(n842) );
  NAND20 U566 ( .A(n859), .B(n122), .Q(n120) );
  NOR21 U567 ( .A(n61), .B(n70), .Q(n59) );
  NAND20 U568 ( .A(n860), .B(n156), .Q(n19) );
  NAND20 U569 ( .A(n839), .B(n71), .Q(n10) );
  INV0 U570 ( .A(n144), .Q(n854) );
  INV0 U571 ( .A(n106), .Q(n848) );
  AOI210 U572 ( .A(n880), .B(n878), .C(n879), .Q(n262) );
  NAND20 U573 ( .A(n895), .B(n224), .Q(n27) );
  INV0 U574 ( .A(n271), .Q(n888) );
  NOR22 U575 ( .A(B[17]), .B(A[17]), .Q(n173) );
  INV1 U576 ( .A(n175), .Q(n865) );
  AOI210 U577 ( .A(n880), .B(n258), .C(n259), .Q(n257) );
  CLKIN3 U578 ( .A(n60), .Q(n838) );
  AOI212 U579 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  INV0 U580 ( .A(n809), .Q(n860) );
  NOR22 U581 ( .A(n809), .B(n162), .Q(n153) );
  INV0 U582 ( .A(n70), .Q(n839) );
  NAND21 U583 ( .A(n836), .B(n62), .Q(n9) );
  NAND20 U584 ( .A(n874), .B(n245), .Q(n30) );
  INV0 U585 ( .A(n244), .Q(n874) );
  AOI210 U586 ( .A(n60), .B(n835), .C(n834), .Q(n47) );
  INV0 U587 ( .A(n260), .Q(n891) );
  NAND20 U588 ( .A(n881), .B(n275), .Q(n36) );
  NAND20 U589 ( .A(n878), .B(n266), .Q(n34) );
  INV0 U590 ( .A(n828), .Q(n895) );
  INV0 U591 ( .A(n231), .Q(n872) );
  INV0 U592 ( .A(n252), .Q(n887) );
  NAND20 U593 ( .A(n887), .B(n253), .Q(n31) );
  NAND20 U594 ( .A(n896), .B(n213), .Q(n26) );
  NAND20 U595 ( .A(n869), .B(n231), .Q(n28) );
  INV0 U596 ( .A(n265), .Q(n878) );
  NAND20 U597 ( .A(n272), .B(n888), .Q(n35) );
  INV0 U598 ( .A(n266), .Q(n879) );
  NAND20 U599 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NOR21 U600 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR22 U601 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NAND20 U602 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U603 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U604 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U605 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND20 U606 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U607 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR20 U608 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NOR20 U609 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U610 ( .A(n111), .B(n55), .Q(n53) );
  NAND20 U611 ( .A(n111), .B(n44), .Q(n42) );
  NOR20 U612 ( .A(n46), .B(n6), .Q(n44) );
  NAND21 U613 ( .A(n175), .B(n21), .Q(n665) );
  NAND22 U614 ( .A(n861), .B(n865), .Q(n666) );
  INV3 U615 ( .A(n21), .Q(n861) );
  NAND22 U616 ( .A(n859), .B(n854), .Q(n140) );
  INV3 U617 ( .A(n59), .Q(n837) );
  INV3 U618 ( .A(n277), .Q(n884) );
  NAND20 U619 ( .A(n866), .B(n177), .Q(n22) );
  NAND22 U620 ( .A(n849), .B(n118), .Q(n15) );
  INV3 U621 ( .A(n832), .Q(n849) );
  NAND22 U622 ( .A(n840), .B(n80), .Q(n11) );
  INV3 U623 ( .A(n79), .Q(n840) );
  NAND22 U624 ( .A(n890), .B(n138), .Q(n17) );
  XOR21 U625 ( .A(n32), .B(n257), .Q(SUM[6]) );
  INV3 U626 ( .A(n255), .Q(n876) );
  XOR20 U627 ( .A(n30), .B(n877), .Q(SUM[8]) );
  NAND22 U628 ( .A(n858), .B(n163), .Q(n20) );
  INV0 U629 ( .A(n172), .Q(n862) );
  INV3 U630 ( .A(n126), .Q(n851) );
  XNR21 U631 ( .A(n34), .B(n880), .Q(SUM[4]) );
  NAND20 U632 ( .A(n893), .B(n206), .Q(n25) );
  XNR21 U633 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND22 U634 ( .A(n843), .B(n89), .Q(n12) );
  INV3 U635 ( .A(n88), .Q(n843) );
  INV3 U636 ( .A(n61), .Q(n836) );
  XNR21 U637 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND22 U638 ( .A(n835), .B(n51), .Q(n8) );
  XNR21 U639 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND22 U640 ( .A(n867), .B(n195), .Q(n24) );
  NAND20 U641 ( .A(n885), .B(n186), .Q(n23) );
  XOR21 U642 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U643 ( .A(n889), .B(n279), .Q(n37) );
  INV3 U644 ( .A(n278), .Q(n889) );
  INV3 U645 ( .A(n99), .Q(n844) );
  XNR21 U646 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NOR21 U647 ( .A(n117), .B(n126), .Q(n115) );
  XOR21 U648 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NOR21 U649 ( .A(n126), .B(n855), .Q(n122) );
  NOR21 U650 ( .A(n88), .B(n845), .Q(n84) );
  NOR21 U651 ( .A(n70), .B(n6), .Q(n66) );
  INV3 U652 ( .A(n107), .Q(n847) );
  AOI210 U653 ( .A(n815), .B(n44), .C(n45), .Q(n43) );
  INV3 U654 ( .A(n51), .Q(n834) );
  AOI210 U655 ( .A(n172), .B(n858), .C(n856), .Q(n159) );
  INV3 U657 ( .A(n163), .Q(n856) );
  AOI211 U658 ( .A(n857), .B(n854), .C(n852), .Q(n141) );
  INV3 U660 ( .A(n145), .Q(n852) );
  INV1 U661 ( .A(n136), .Q(n853) );
  XOR21 U662 ( .A(n36), .B(n884), .Q(SUM[2]) );
  INV3 U663 ( .A(n274), .Q(n881) );
  XNR21 U664 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NOR21 U666 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR21 U667 ( .A(B[28]), .B(A[28]), .Q(n70) );
  XNR21 U668 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U669 ( .A(n833), .B(n40), .Q(n7) );
  NOR21 U670 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND22 U671 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U672 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U673 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NOR20 U674 ( .A(B[2]), .B(A[2]), .Q(n274) );
  INV3 U675 ( .A(n39), .Q(n833) );
  INV3 U676 ( .A(n50), .Q(n835) );
  INV3 U677 ( .A(n38), .Q(SUM[0]) );
  NAND22 U678 ( .A(n883), .B(n281), .Q(n38) );
  INV3 U679 ( .A(n280), .Q(n883) );
  NOR20 U680 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U681 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U682 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND22 U683 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NOR20 U684 ( .A(B[1]), .B(A[1]), .Q(n278) );
  AOI210 U685 ( .A(n871), .B(n203), .C(n830), .Q(n198) );
  INV1 U686 ( .A(n811), .Q(n880) );
endmodule


module adder_26 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_26_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_25_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n52, n53, n54, n57, n58, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n79, n80, n81, n82, n83, n84, n85, n88,
         n89, n90, n93, n94, n99, n100, n101, n102, n103, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n121, n122, n123, n124, n125, n126, n131, n132, n133, n134, n135,
         n138, n139, n140, n141, n142, n147, n148, n149, n150, n151, n152,
         n153, n156, n157, n158, n161, n162, n167, n168, n169, n170, n171,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n186, n187, n188, n189, n194, n195, n196, n199, n200, n202, n203,
         n204, n205, n206, n207, n208, n209, n212, n213, n214, n215, n216,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n240, n241, n243, n244, n245, n246,
         n247, n248, n249, n250, n252, n253, n254, n255, n256, n397, n737,
         n738, n739, n740, n741, n742, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807;

  OAI212 U16 ( .A(n53), .B(n45), .C(n46), .Q(n44) );
  OAI212 U40 ( .A(n71), .B(n63), .C(n64), .Q(n62) );
  OAI212 U46 ( .A(n66), .B(n742), .C(n67), .Q(n65) );
  OAI212 U70 ( .A(n84), .B(n742), .C(n85), .Q(n83) );
  OAI212 U80 ( .A(n801), .B(n742), .C(n799), .Q(n90) );
  OAI212 U102 ( .A(n142), .B(n107), .C(n108), .Q(n106) );
  AOI212 U154 ( .A(n147), .B(n162), .C(n148), .Q(n142) );
  OAI212 U180 ( .A(n171), .B(n167), .C(n168), .Q(n162) );
  OAI212 U193 ( .A(n174), .B(n202), .C(n175), .Q(n173) );
  OAI212 U219 ( .A(n200), .B(n194), .C(n195), .Q(n189) );
  OAI212 U236 ( .A(n209), .B(n205), .C(n206), .Q(n204) );
  OAI212 U242 ( .A(n208), .B(n747), .C(n209), .Q(n207) );
  OAI212 U252 ( .A(n215), .B(n747), .C(n216), .Q(n214) );
  OAI212 U263 ( .A(n223), .B(n243), .C(n224), .Q(n222) );
  OAI212 U267 ( .A(n231), .B(n227), .C(n228), .Q(n226) );
  OAI212 U273 ( .A(n230), .B(n232), .C(n231), .Q(n229) );
  OAI212 U281 ( .A(n241), .B(n235), .C(n236), .Q(n234) );
  OAI212 U298 ( .A(n250), .B(n246), .C(n247), .Q(n245) );
  OAI212 U304 ( .A(n249), .B(n745), .C(n250), .Q(n248) );
  OAI212 U311 ( .A(n256), .B(n253), .C(n254), .Q(n252) );
  OAI212 U387 ( .A(n114), .B(n749), .C(n115), .Q(n113) );
  AOI212 U398 ( .A(n173), .B(n105), .C(n106), .Q(n1) );
  OAI212 U349 ( .A(n774), .B(n74), .C(n771), .Q(n58) );
  OAI212 U358 ( .A(n773), .B(n742), .C(n770), .Q(n54) );
  OAI212 U392 ( .A(n103), .B(n99), .C(n100), .Q(n94) );
  OAI212 U406 ( .A(n131), .B(n139), .C(n132), .Q(n126) );
  AOI212 U337 ( .A(n94), .B(n79), .C(n80), .Q(n74) );
  OAI212 U354 ( .A(n765), .B(n742), .C(n766), .Q(n36) );
  OAI212 U410 ( .A(n788), .B(n749), .C(n789), .Q(n158) );
  AOI212 U325 ( .A(n189), .B(n176), .C(n177), .Q(n175) );
  OAI212 U386 ( .A(n89), .B(n741), .C(n82), .Q(n80) );
  OAI212 U412 ( .A(n102), .B(n742), .C(n103), .Q(n101) );
  OAI212 U370 ( .A(n152), .B(n749), .C(n153), .Q(n151) );
  XNR22 U324 ( .A(n16), .B(n158), .Q(SUM[17]) );
  XOR22 U326 ( .A(n19), .B(n180), .Q(SUM[14]) );
  NOR24 U327 ( .A(n178), .B(n183), .Q(n176) );
  NOR23 U328 ( .A(B[13]), .B(A[13]), .Q(n183) );
  XOR22 U329 ( .A(n10), .B(n742), .Q(SUM[23]) );
  NOR24 U330 ( .A(B[12]), .B(A[12]), .Q(n194) );
  NAND23 U331 ( .A(n161), .B(n147), .Q(n141) );
  NOR22 U332 ( .A(n167), .B(n170), .Q(n161) );
  OAI211 U333 ( .A(n749), .B(n123), .C(n124), .Q(n122) );
  XNR22 U334 ( .A(n13), .B(n133), .Q(SUM[20]) );
  NOR23 U335 ( .A(A[14]), .B(B[14]), .Q(n178) );
  NOR23 U336 ( .A(B[16]), .B(A[16]), .Q(n167) );
  NOR22 U338 ( .A(B[15]), .B(A[15]), .Q(n170) );
  NOR22 U339 ( .A(n111), .B(n118), .Q(n109) );
  NOR22 U340 ( .A(n131), .B(n138), .Q(n125) );
  NOR22 U341 ( .A(n149), .B(n156), .Q(n147) );
  NAND22 U342 ( .A(A[11]), .B(B[11]), .Q(n200) );
  XOR21 U343 ( .A(n18), .B(n749), .Q(SUM[15]) );
  NOR22 U344 ( .A(B[22]), .B(A[22]), .Q(n111) );
  NAND20 U345 ( .A(B[20]), .B(A[20]), .Q(n132) );
  NOR22 U346 ( .A(B[20]), .B(A[20]), .Q(n131) );
  NOR22 U347 ( .A(B[21]), .B(A[21]), .Q(n118) );
  NOR22 U348 ( .A(n107), .B(n141), .Q(n105) );
  NAND22 U350 ( .A(n8), .B(n90), .Q(n739) );
  NAND26 U351 ( .A(n737), .B(n738), .Q(n740) );
  NAND28 U352 ( .A(n739), .B(n740), .Q(SUM[25]) );
  INV6 U353 ( .A(n8), .Q(n737) );
  CLKIN6 U355 ( .A(n90), .Q(n738) );
  NAND22 U356 ( .A(n791), .B(n89), .Q(n8) );
  INV0 U357 ( .A(n183), .Q(n779) );
  OAI210 U359 ( .A(n183), .B(n793), .C(n186), .Q(n182) );
  NAND24 U360 ( .A(n397), .B(n150), .Q(n148) );
  INV0 U361 ( .A(n111), .Q(n796) );
  NOR20 U362 ( .A(B[27]), .B(A[27]), .Q(n70) );
  NAND21 U363 ( .A(A[12]), .B(B[12]), .Q(n195) );
  NOR20 U364 ( .A(B[11]), .B(A[11]), .Q(n199) );
  OAI212 U365 ( .A(n48), .B(n742), .C(n49), .Q(n47) );
  BUF15 U366 ( .A(n1), .Q(n742) );
  XNR22 U367 ( .A(n3), .B(n47), .Q(SUM[30]) );
  AOI211 U368 ( .A(n58), .B(n768), .C(n767), .Q(n49) );
  XNR22 U369 ( .A(n11), .B(n113), .Q(SUM[22]) );
  NAND20 U371 ( .A(n782), .B(n139), .Q(n14) );
  INV0 U372 ( .A(n139), .Q(n780) );
  NAND20 U373 ( .A(B[22]), .B(A[22]), .Q(n112) );
  NOR22 U374 ( .A(B[23]), .B(A[23]), .Q(n102) );
  OAI212 U375 ( .A(n186), .B(n178), .C(n179), .Q(n177) );
  NAND22 U376 ( .A(A[13]), .B(B[13]), .Q(n186) );
  NAND22 U377 ( .A(B[18]), .B(A[18]), .Q(n150) );
  XNR22 U378 ( .A(n4), .B(n54), .Q(SUM[29]) );
  NAND21 U379 ( .A(A[25]), .B(B[25]), .Q(n89) );
  NOR22 U380 ( .A(n741), .B(n88), .Q(n79) );
  NAND22 U381 ( .A(A[15]), .B(B[15]), .Q(n171) );
  NAND22 U382 ( .A(n57), .B(n768), .Q(n48) );
  NAND20 U383 ( .A(n805), .B(n132), .Q(n13) );
  OAI212 U384 ( .A(n73), .B(n742), .C(n74), .Q(n72) );
  OAI211 U385 ( .A(n118), .B(n781), .C(n121), .Q(n117) );
  INV0 U388 ( .A(n118), .Q(n797) );
  NOR21 U389 ( .A(n118), .B(n783), .Q(n116) );
  XNR22 U390 ( .A(n6), .B(n72), .Q(SUM[27]) );
  NAND21 U391 ( .A(A[21]), .B(B[21]), .Q(n121) );
  CLKIN6 U393 ( .A(n149), .Q(n785) );
  NOR22 U394 ( .A(B[18]), .B(A[18]), .Q(n149) );
  NOR22 U395 ( .A(B[17]), .B(A[17]), .Q(n156) );
  XNR22 U396 ( .A(n14), .B(n140), .Q(SUM[19]) );
  NAND21 U397 ( .A(n787), .B(n171), .Q(n18) );
  OAI211 U399 ( .A(n170), .B(n749), .C(n171), .Q(n169) );
  NAND21 U400 ( .A(A[14]), .B(B[14]), .Q(n179) );
  OAI211 U401 ( .A(n121), .B(n111), .C(n112), .Q(n110) );
  NAND22 U402 ( .A(A[16]), .B(B[16]), .Q(n168) );
  XNR22 U403 ( .A(n7), .B(n83), .Q(SUM[26]) );
  AOI211 U404 ( .A(n126), .B(n109), .C(n110), .Q(n108) );
  XNR22 U405 ( .A(n5), .B(n65), .Q(SUM[28]) );
  XNR22 U407 ( .A(n9), .B(n101), .Q(SUM[24]) );
  NAND22 U408 ( .A(A[17]), .B(B[17]), .Q(n157) );
  INV0 U409 ( .A(n167), .Q(n802) );
  INV0 U411 ( .A(n131), .Q(n805) );
  NAND21 U413 ( .A(n786), .B(n116), .Q(n114) );
  INV3 U414 ( .A(n141), .Q(n786) );
  OAI211 U415 ( .A(n134), .B(n749), .C(n135), .Q(n133) );
  BUF6 U416 ( .A(n81), .Q(n741) );
  INV0 U417 ( .A(n138), .Q(n782) );
  NAND21 U418 ( .A(A[19]), .B(B[19]), .Q(n139) );
  INV0 U419 ( .A(n73), .Q(n776) );
  NAND20 U420 ( .A(n786), .B(n782), .Q(n134) );
  INV1 U421 ( .A(n71), .Q(n769) );
  NAND20 U422 ( .A(n807), .B(n64), .Q(n5) );
  INV1 U423 ( .A(n70), .Q(n772) );
  AOI210 U424 ( .A(n784), .B(n782), .C(n780), .Q(n135) );
  NAND20 U425 ( .A(n786), .B(n125), .Q(n123) );
  NAND20 U426 ( .A(n93), .B(n791), .Q(n84) );
  NAND20 U427 ( .A(n797), .B(n121), .Q(n12) );
  NAND20 U428 ( .A(A[4]), .B(B[4]), .Q(n241) );
  NAND20 U429 ( .A(A[8]), .B(B[8]), .Q(n216) );
  NAND20 U430 ( .A(A[9]), .B(B[9]), .Q(n213) );
  NOR20 U431 ( .A(n41), .B(n73), .Q(n39) );
  CLKIN3 U432 ( .A(n58), .Q(n770) );
  CLKIN0 U433 ( .A(n161), .Q(n788) );
  NOR21 U434 ( .A(n99), .B(n102), .Q(n93) );
  NAND20 U435 ( .A(n188), .B(n176), .Q(n174) );
  INV3 U436 ( .A(n74), .Q(n777) );
  NAND20 U437 ( .A(n161), .B(n804), .Q(n152) );
  NAND20 U438 ( .A(n785), .B(n150), .Q(n15) );
  NAND20 U439 ( .A(n794), .B(n200), .Q(n22) );
  INV0 U440 ( .A(n194), .Q(n798) );
  INV0 U441 ( .A(n178), .Q(n778) );
  INV0 U442 ( .A(n170), .Q(n787) );
  INV0 U443 ( .A(n53), .Q(n767) );
  INV3 U444 ( .A(n52), .Q(n768) );
  NOR21 U445 ( .A(n63), .B(n70), .Q(n61) );
  INV0 U446 ( .A(n200), .Q(n792) );
  NOR20 U447 ( .A(B[26]), .B(A[26]), .Q(n81) );
  NAND20 U448 ( .A(A[27]), .B(B[27]), .Q(n71) );
  NOR20 U449 ( .A(B[30]), .B(A[30]), .Q(n45) );
  NOR20 U450 ( .A(B[10]), .B(A[10]), .Q(n205) );
  NAND20 U451 ( .A(A[26]), .B(B[26]), .Q(n82) );
  NAND20 U452 ( .A(B[31]), .B(A[31]), .Q(n35) );
  NOR21 U453 ( .A(n774), .B(n73), .Q(n57) );
  INV3 U454 ( .A(n39), .Q(n765) );
  INV3 U455 ( .A(n62), .Q(n771) );
  NAND22 U456 ( .A(n93), .B(n79), .Q(n73) );
  AOI211 U457 ( .A(n784), .B(n125), .C(n126), .Q(n124) );
  INV6 U458 ( .A(n173), .Q(n749) );
  NAND22 U459 ( .A(n61), .B(n43), .Q(n41) );
  NAND22 U460 ( .A(n125), .B(n109), .Q(n107) );
  CLKIN2 U461 ( .A(n142), .Q(n784) );
  INV3 U462 ( .A(n61), .Q(n774) );
  INV3 U463 ( .A(n93), .Q(n801) );
  NAND22 U464 ( .A(n776), .B(n772), .Q(n66) );
  AOI211 U465 ( .A(n746), .B(n233), .C(n234), .Q(n232) );
  INV3 U466 ( .A(n222), .Q(n747) );
  INV3 U467 ( .A(n202), .Q(n748) );
  INV3 U468 ( .A(n243), .Q(n746) );
  INV3 U469 ( .A(n252), .Q(n745) );
  XOR21 U470 ( .A(n20), .B(n187), .Q(SUM[13]) );
  NAND22 U471 ( .A(n779), .B(n186), .Q(n20) );
  NAND22 U472 ( .A(n803), .B(n785), .Q(n397) );
  NAND22 U473 ( .A(n768), .B(n53), .Q(n4) );
  CLKIN3 U474 ( .A(n57), .Q(n773) );
  XNR21 U475 ( .A(n17), .B(n169), .Q(SUM[16]) );
  NAND22 U476 ( .A(n802), .B(n168), .Q(n17) );
  NAND22 U477 ( .A(n804), .B(n157), .Q(n16) );
  INV0 U478 ( .A(n162), .Q(n789) );
  NAND20 U479 ( .A(n796), .B(n112), .Q(n11) );
  XNR21 U480 ( .A(n15), .B(n151), .Q(SUM[18]) );
  NAND22 U481 ( .A(n775), .B(n82), .Q(n7) );
  INV3 U482 ( .A(n741), .Q(n775) );
  INV0 U483 ( .A(n63), .Q(n807) );
  NAND22 U484 ( .A(n764), .B(n46), .Q(n3) );
  INV3 U485 ( .A(n45), .Q(n764) );
  XNR21 U486 ( .A(n23), .B(n207), .Q(SUM[10]) );
  NAND22 U487 ( .A(n762), .B(n206), .Q(n23) );
  INV3 U488 ( .A(n205), .Q(n762) );
  NOR21 U489 ( .A(n45), .B(n52), .Q(n43) );
  NAND20 U490 ( .A(n806), .B(n103), .Q(n10) );
  INV2 U491 ( .A(n102), .Q(n806) );
  NAND22 U492 ( .A(n772), .B(n71), .Q(n6) );
  NAND20 U493 ( .A(n800), .B(n100), .Q(n9) );
  INV0 U494 ( .A(n99), .Q(n800) );
  XNR21 U495 ( .A(n12), .B(n122), .Q(SUM[21]) );
  XNR21 U496 ( .A(n22), .B(n748), .Q(SUM[11]) );
  CLKIN0 U497 ( .A(n94), .Q(n799) );
  INV2 U498 ( .A(n125), .Q(n783) );
  INV0 U499 ( .A(n189), .Q(n793) );
  NAND22 U500 ( .A(n778), .B(n179), .Q(n19) );
  AOI211 U501 ( .A(n748), .B(n181), .C(n182), .Q(n180) );
  XOR21 U502 ( .A(n21), .B(n196), .Q(SUM[12]) );
  NAND20 U503 ( .A(n195), .B(n798), .Q(n21) );
  AOI211 U504 ( .A(n748), .B(n794), .C(n792), .Q(n196) );
  CLKIN1 U505 ( .A(n88), .Q(n791) );
  AOI210 U506 ( .A(n94), .B(n791), .C(n790), .Q(n85) );
  INV3 U507 ( .A(n89), .Q(n790) );
  AOI210 U508 ( .A(n784), .B(n116), .C(n117), .Q(n115) );
  CLKIN0 U509 ( .A(n126), .Q(n781) );
  CLKIN3 U510 ( .A(n199), .Q(n794) );
  CLKIN2 U511 ( .A(n40), .Q(n766) );
  AOI210 U512 ( .A(n62), .B(n43), .C(n44), .Q(n42) );
  INV3 U513 ( .A(n156), .Q(n804) );
  AOI211 U514 ( .A(n777), .B(n772), .C(n769), .Q(n67) );
  INV3 U515 ( .A(n157), .Q(n803) );
  XOR21 U516 ( .A(n28), .B(n237), .Q(SUM[5]) );
  NAND22 U517 ( .A(n755), .B(n236), .Q(n28) );
  AOI211 U518 ( .A(n746), .B(n754), .C(n753), .Q(n237) );
  INV3 U519 ( .A(n235), .Q(n755) );
  XOR21 U520 ( .A(n31), .B(n745), .Q(SUM[2]) );
  NAND22 U521 ( .A(n751), .B(n250), .Q(n31) );
  INV3 U522 ( .A(n249), .Q(n751) );
  XOR21 U523 ( .A(n27), .B(n232), .Q(SUM[6]) );
  NAND22 U524 ( .A(n756), .B(n231), .Q(n27) );
  INV3 U525 ( .A(n230), .Q(n756) );
  XOR21 U526 ( .A(n25), .B(n747), .Q(SUM[8]) );
  NAND22 U527 ( .A(n759), .B(n216), .Q(n25) );
  XOR21 U528 ( .A(n256), .B(n32), .Q(SUM[1]) );
  NAND22 U529 ( .A(n750), .B(n254), .Q(n32) );
  INV3 U530 ( .A(n253), .Q(n750) );
  NAND22 U531 ( .A(n233), .B(n225), .Q(n223) );
  AOI211 U532 ( .A(n234), .B(n225), .C(n226), .Q(n224) );
  NOR21 U533 ( .A(n227), .B(n230), .Q(n225) );
  AOI211 U534 ( .A(n203), .B(n222), .C(n204), .Q(n202) );
  NOR21 U535 ( .A(n208), .B(n205), .Q(n203) );
  XNR21 U536 ( .A(n26), .B(n229), .Q(SUM[7]) );
  NAND22 U537 ( .A(n757), .B(n228), .Q(n26) );
  INV3 U538 ( .A(n227), .Q(n757) );
  XNR21 U539 ( .A(n30), .B(n248), .Q(SUM[3]) );
  NAND22 U540 ( .A(n752), .B(n247), .Q(n30) );
  INV3 U541 ( .A(n246), .Q(n752) );
  XNR21 U542 ( .A(n24), .B(n214), .Q(SUM[9]) );
  NAND22 U543 ( .A(n761), .B(n213), .Q(n24) );
  AOI211 U544 ( .A(n252), .B(n244), .C(n245), .Q(n243) );
  NOR21 U545 ( .A(n246), .B(n249), .Q(n244) );
  XNR21 U546 ( .A(n29), .B(n746), .Q(SUM[4]) );
  NAND22 U547 ( .A(n754), .B(n241), .Q(n29) );
  NOR20 U548 ( .A(n194), .B(n199), .Q(n188) );
  AOI211 U549 ( .A(n761), .B(n758), .C(n760), .Q(n209) );
  INV3 U550 ( .A(n216), .Q(n758) );
  INV3 U551 ( .A(n213), .Q(n760) );
  NOR21 U552 ( .A(n235), .B(n240), .Q(n233) );
  NOR21 U553 ( .A(n183), .B(n795), .Q(n181) );
  INV3 U554 ( .A(n188), .Q(n795) );
  NAND22 U555 ( .A(n759), .B(n761), .Q(n208) );
  INV3 U556 ( .A(n215), .Q(n759) );
  INV3 U557 ( .A(n240), .Q(n754) );
  INV3 U558 ( .A(n241), .Q(n753) );
  XNR21 U559 ( .A(n2), .B(n36), .Q(SUM[31]) );
  NAND22 U560 ( .A(n763), .B(n35), .Q(n2) );
  NAND20 U561 ( .A(A[28]), .B(B[28]), .Q(n64) );
  INV3 U562 ( .A(n34), .Q(n763) );
  NOR20 U563 ( .A(A[31]), .B(B[31]), .Q(n34) );
  NAND20 U564 ( .A(A[10]), .B(B[10]), .Q(n206) );
  INV3 U565 ( .A(n212), .Q(n761) );
  NOR20 U566 ( .A(B[9]), .B(A[9]), .Q(n212) );
  INV3 U567 ( .A(n33), .Q(SUM[0]) );
  NAND22 U568 ( .A(n744), .B(n256), .Q(n33) );
  INV3 U569 ( .A(n255), .Q(n744) );
  NOR20 U570 ( .A(B[0]), .B(A[0]), .Q(n255) );
  NOR20 U571 ( .A(B[3]), .B(A[3]), .Q(n246) );
  NOR20 U572 ( .A(B[7]), .B(A[7]), .Q(n227) );
  NOR20 U573 ( .A(B[5]), .B(A[5]), .Q(n235) );
  NOR20 U574 ( .A(B[2]), .B(A[2]), .Q(n249) );
  NOR20 U575 ( .A(B[6]), .B(A[6]), .Q(n230) );
  NAND20 U576 ( .A(A[0]), .B(B[0]), .Q(n256) );
  NAND20 U577 ( .A(A[2]), .B(B[2]), .Q(n250) );
  NAND20 U578 ( .A(A[6]), .B(B[6]), .Q(n231) );
  NOR20 U579 ( .A(B[4]), .B(A[4]), .Q(n240) );
  NOR20 U580 ( .A(B[1]), .B(A[1]), .Q(n253) );
  NOR20 U581 ( .A(B[8]), .B(A[8]), .Q(n215) );
  NAND20 U582 ( .A(A[1]), .B(B[1]), .Q(n254) );
  NAND20 U583 ( .A(A[3]), .B(B[3]), .Q(n247) );
  NAND20 U584 ( .A(A[5]), .B(B[5]), .Q(n236) );
  NAND20 U585 ( .A(A[7]), .B(B[7]), .Q(n228) );
  NOR20 U586 ( .A(B[29]), .B(A[29]), .Q(n52) );
  NAND21 U587 ( .A(A[29]), .B(B[29]), .Q(n53) );
  NAND21 U588 ( .A(A[30]), .B(B[30]), .Q(n46) );
  NAND21 U589 ( .A(A[23]), .B(B[23]), .Q(n103) );
  OAI210 U590 ( .A(n41), .B(n74), .C(n42), .Q(n40) );
  NOR21 U591 ( .A(B[25]), .B(A[25]), .Q(n88) );
  NAND22 U592 ( .A(A[24]), .B(B[24]), .Q(n100) );
  NOR22 U593 ( .A(A[19]), .B(B[19]), .Q(n138) );
  AOI211 U594 ( .A(n748), .B(n188), .C(n189), .Q(n187) );
  OAI211 U595 ( .A(n141), .B(n749), .C(n142), .Q(n140) );
  AOI210 U596 ( .A(n162), .B(n804), .C(n803), .Q(n153) );
  NOR21 U597 ( .A(B[28]), .B(A[28]), .Q(n63) );
  NOR22 U598 ( .A(B[24]), .B(A[24]), .Q(n99) );
endmodule


module adder_25 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_25_DW01_add_2 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_24_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n416, n422,
         n424, n425, n494, n632, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n834;

  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U391 ( .A(n223), .B(n231), .C(n224), .Q(n222) );
  OAI212 U490 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U493 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  AOI212 U407 ( .A(n98), .B(n77), .C(n78), .Q(n494) );
  OAI212 U410 ( .A(n770), .B(n102), .C(n103), .Q(n101) );
  OAI212 U413 ( .A(n73), .B(n770), .C(n74), .Q(n72) );
  OAI212 U430 ( .A(n770), .B(n82), .C(n83), .Q(n81) );
  OAI212 U438 ( .A(n770), .B(n53), .C(n54), .Q(n52) );
  OAI212 U467 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  AOI212 U508 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U427 ( .A(n176), .B(n770), .C(n177), .Q(n175) );
  OAI212 U428 ( .A(n772), .B(n770), .C(n775), .Q(n164) );
  OAI212 U429 ( .A(n158), .B(n770), .C(n159), .Q(n157) );
  OAI212 U494 ( .A(n129), .B(n770), .C(n130), .Q(n128) );
  OAI212 U450 ( .A(n120), .B(n770), .C(n121), .Q(n119) );
  OAI212 U497 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U483 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U477 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U459 ( .A(n88), .B(n786), .C(n89), .Q(n85) );
  OAI212 U433 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U488 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U398 ( .A(n126), .B(n783), .C(n127), .Q(n123) );
  NAND23 U349 ( .A(n239), .B(n221), .Q(n219) );
  NOR22 U350 ( .A(n241), .B(n244), .Q(n239) );
  INV1 U351 ( .A(n220), .Q(n813) );
  NAND22 U352 ( .A(n258), .B(n250), .Q(n248) );
  NOR22 U353 ( .A(n265), .B(n260), .Q(n258) );
  NOR23 U354 ( .A(n61), .B(n70), .Q(n59) );
  NAND22 U355 ( .A(n111), .B(n66), .Q(n64) );
  AOI212 U356 ( .A(n769), .B(n66), .C(n67), .Q(n65) );
  AOI212 U357 ( .A(n769), .B(n789), .C(n788), .Q(n103) );
  INV3 U358 ( .A(n106), .Q(n789) );
  XNR22 U359 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NOR23 U360 ( .A(B[27]), .B(A[27]), .Q(n79) );
  OAI210 U361 ( .A(n194), .B(n811), .C(n195), .Q(n191) );
  INV6 U362 ( .A(n416), .Q(n822) );
  INV3 U363 ( .A(n203), .Q(n809) );
  AOI212 U364 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NAND26 U365 ( .A(n97), .B(n77), .Q(n6) );
  NAND22 U366 ( .A(n111), .B(n97), .Q(n91) );
  NOR23 U367 ( .A(n99), .B(n106), .Q(n97) );
  NAND28 U368 ( .A(n203), .B(n183), .Q(n181) );
  NOR24 U369 ( .A(n181), .B(n219), .Q(n179) );
  NOR23 U370 ( .A(n205), .B(n212), .Q(n203) );
  NOR22 U371 ( .A(n173), .B(n176), .Q(n171) );
  AOI212 U372 ( .A(n172), .B(n153), .C(n632), .Q(n425) );
  NAND24 U373 ( .A(n422), .B(n174), .Q(n172) );
  OAI212 U374 ( .A(n163), .B(n155), .C(n156), .Q(n632) );
  NOR22 U375 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR23 U376 ( .A(n137), .B(n144), .Q(n135) );
  NOR22 U377 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR23 U378 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR24 U379 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND24 U380 ( .A(n171), .B(n153), .Q(n151) );
  NOR24 U381 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NAND22 U382 ( .A(n773), .B(n135), .Q(n129) );
  INV1 U383 ( .A(n151), .Q(n773) );
  NAND24 U384 ( .A(n135), .B(n115), .Q(n113) );
  NOR24 U385 ( .A(n117), .B(n126), .Q(n115) );
  NOR24 U386 ( .A(n79), .B(n88), .Q(n77) );
  INV2 U387 ( .A(n98), .Q(n786) );
  NOR23 U388 ( .A(n252), .B(n255), .Q(n250) );
  NOR22 U389 ( .A(n88), .B(n790), .Q(n84) );
  NOR22 U390 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR21 U392 ( .A(n70), .B(n6), .Q(n66) );
  INV3 U393 ( .A(n59), .Q(n794) );
  NOR23 U394 ( .A(B[22]), .B(A[22]), .Q(n126) );
  INV3 U395 ( .A(n425), .Q(n776) );
  INV3 U396 ( .A(n97), .Q(n790) );
  NAND24 U397 ( .A(n424), .B(n100), .Q(n98) );
  NOR23 U399 ( .A(n113), .B(n151), .Q(n111) );
  NOR23 U400 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NOR22 U401 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR22 U402 ( .A(B[14]), .B(A[14]), .Q(n194) );
  INV3 U403 ( .A(n50), .Q(n800) );
  NOR21 U404 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U405 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND22 U406 ( .A(A[26]), .B(B[26]), .Q(n89) );
  INV3 U408 ( .A(n268), .Q(n828) );
  NAND22 U409 ( .A(B[6]), .B(A[6]), .Q(n256) );
  NAND22 U411 ( .A(A[16]), .B(B[16]), .Q(n177) );
  AOI212 U412 ( .A(n769), .B(n44), .C(n45), .Q(n43) );
  INV2 U414 ( .A(n775), .Q(n768) );
  CLKIN1 U415 ( .A(n172), .Q(n775) );
  NOR23 U416 ( .A(A[17]), .B(B[17]), .Q(n173) );
  NAND22 U417 ( .A(A[19]), .B(B[19]), .Q(n156) );
  AOI212 U418 ( .A(n769), .B(n791), .C(n787), .Q(n74) );
  NAND24 U419 ( .A(n778), .B(n805), .Q(n422) );
  XNR22 U420 ( .A(n7), .B(n41), .Q(SUM[31]) );
  XNR22 U421 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XOR21 U422 ( .A(n22), .B(n770), .Q(SUM[16]) );
  XNR22 U423 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND21 U424 ( .A(n800), .B(n51), .Q(n8) );
  XOR20 U425 ( .A(n30), .B(n822), .Q(SUM[8]) );
  OAI211 U426 ( .A(n244), .B(n822), .C(n245), .Q(n243) );
  OAI211 U431 ( .A(n188), .B(n822), .C(n189), .Q(n187) );
  OAI211 U432 ( .A(n208), .B(n822), .C(n209), .Q(n207) );
  OAI211 U434 ( .A(n197), .B(n822), .C(n198), .Q(n196) );
  OAI211 U435 ( .A(n820), .B(n822), .C(n818), .Q(n232) );
  OAI211 U436 ( .A(n226), .B(n822), .C(n227), .Q(n225) );
  NAND21 U437 ( .A(A[4]), .B(B[4]), .Q(n266) );
  OAI211 U439 ( .A(n219), .B(n822), .C(n220), .Q(n214) );
  BUF15 U440 ( .A(n112), .Q(n769) );
  AOI212 U441 ( .A(n769), .B(n97), .C(n98), .Q(n92) );
  XNR22 U442 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NAND21 U443 ( .A(A[23]), .B(B[23]), .Q(n118) );
  OAI212 U444 ( .A(n494), .B(n46), .C(n47), .Q(n45) );
  NAND22 U445 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND21 U446 ( .A(A[13]), .B(B[13]), .Q(n206) );
  OAI212 U447 ( .A(n794), .B(n5), .C(n795), .Q(n56) );
  NAND21 U448 ( .A(n773), .B(n803), .Q(n140) );
  NAND21 U449 ( .A(A[29]), .B(B[29]), .Q(n62) );
  OAI212 U451 ( .A(n140), .B(n770), .C(n141), .Q(n139) );
  NAND21 U452 ( .A(n803), .B(n145), .Q(n18) );
  NAND22 U453 ( .A(B[20]), .B(A[20]), .Q(n145) );
  NAND22 U454 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND21 U455 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND24 U456 ( .A(n59), .B(n800), .Q(n46) );
  OAI212 U457 ( .A(n151), .B(n770), .C(n425), .Q(n146) );
  NAND21 U458 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND22 U460 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NOR23 U461 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NAND22 U462 ( .A(n111), .B(n55), .Q(n53) );
  NOR22 U463 ( .A(n794), .B(n6), .Q(n55) );
  NOR22 U464 ( .A(n126), .B(n782), .Q(n122) );
  CLKIN3 U465 ( .A(n135), .Q(n782) );
  NAND21 U466 ( .A(n773), .B(n122), .Q(n120) );
  NOR24 U468 ( .A(A[25]), .B(B[25]), .Q(n99) );
  XNR22 U469 ( .A(n9), .B(n63), .Q(SUM[29]) );
  OAI212 U470 ( .A(n64), .B(n770), .C(n65), .Q(n63) );
  NOR24 U471 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND21 U472 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND21 U473 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND22 U474 ( .A(A[10]), .B(B[10]), .Q(n231) );
  AOI210 U475 ( .A(n776), .B(n135), .C(n136), .Q(n130) );
  CLKIN3 U476 ( .A(n145), .Q(n802) );
  NOR22 U478 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NAND21 U479 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NOR24 U480 ( .A(n155), .B(n162), .Q(n153) );
  NOR22 U481 ( .A(B[18]), .B(A[18]), .Q(n162) );
  CLKBU15 U482 ( .A(n178), .Q(n770) );
  NOR24 U484 ( .A(B[19]), .B(A[19]), .Q(n155) );
  INV1 U485 ( .A(n155), .Q(n804) );
  NAND21 U486 ( .A(A[21]), .B(B[21]), .Q(n138) );
  CLKIN1 U487 ( .A(n136), .Q(n783) );
  OAI212 U489 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  NAND22 U491 ( .A(A[28]), .B(B[28]), .Q(n71) );
  INV1 U492 ( .A(n162), .Q(n779) );
  OAI212 U495 ( .A(n774), .B(n770), .C(n777), .Q(n108) );
  INV1 U496 ( .A(n111), .Q(n774) );
  NAND22 U498 ( .A(n111), .B(n44), .Q(n42) );
  NOR22 U499 ( .A(n46), .B(n6), .Q(n44) );
  OAI211 U500 ( .A(n248), .B(n268), .C(n249), .Q(n416) );
  AOI212 U501 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U502 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  NOR23 U503 ( .A(n223), .B(n230), .Q(n221) );
  INV0 U504 ( .A(n223), .Q(n814) );
  NAND21 U505 ( .A(B[25]), .B(A[25]), .Q(n100) );
  OAI212 U506 ( .A(n91), .B(n770), .C(n92), .Q(n90) );
  NAND21 U507 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV0 U509 ( .A(n213), .Q(n810) );
  CLKIN1 U510 ( .A(n204), .Q(n811) );
  NAND21 U511 ( .A(n111), .B(n789), .Q(n102) );
  AOI212 U512 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  NAND21 U513 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NOR24 U514 ( .A(n185), .B(n194), .Q(n183) );
  OAI212 U515 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  NAND21 U516 ( .A(n111), .B(n84), .Q(n82) );
  INV2 U517 ( .A(n6), .Q(n791) );
  NAND22 U518 ( .A(n111), .B(n791), .Q(n73) );
  OAI210 U519 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  AOI211 U520 ( .A(n828), .B(n258), .C(n259), .Q(n257) );
  OAI212 U521 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  AOI212 U522 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  AOI212 U523 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  AOI210 U524 ( .A(n768), .B(n779), .C(n780), .Q(n159) );
  AOI211 U525 ( .A(n769), .B(n84), .C(n85), .Q(n83) );
  OAI212 U526 ( .A(n42), .B(n770), .C(n43), .Q(n41) );
  NAND22 U527 ( .A(n815), .B(n203), .Q(n197) );
  CLKIN6 U528 ( .A(n173), .Q(n805) );
  NOR22 U529 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NAND22 U530 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NOR22 U531 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR22 U532 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR22 U533 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NAND22 U534 ( .A(A[1]), .B(B[1]), .Q(n279) );
  INV0 U535 ( .A(n171), .Q(n772) );
  INV3 U536 ( .A(n494), .Q(n787) );
  INV0 U537 ( .A(n239), .Q(n820) );
  CLKIN1 U538 ( .A(n60), .Q(n795) );
  INV0 U539 ( .A(n144), .Q(n803) );
  NAND22 U540 ( .A(n815), .B(n190), .Q(n188) );
  INV0 U541 ( .A(n277), .Q(n832) );
  INV0 U542 ( .A(n278), .Q(n831) );
  AOI210 U543 ( .A(n813), .B(n203), .C(n204), .Q(n198) );
  AOI211 U544 ( .A(n813), .B(n190), .C(n191), .Q(n189) );
  AOI210 U545 ( .A(n828), .B(n826), .C(n827), .Q(n262) );
  INV0 U546 ( .A(n266), .Q(n827) );
  OAI210 U547 ( .A(n274), .B(n832), .C(n275), .Q(n273) );
  INV0 U548 ( .A(n230), .Q(n816) );
  INV0 U549 ( .A(n265), .Q(n826) );
  INV0 U550 ( .A(n274), .Q(n829) );
  INV0 U551 ( .A(n271), .Q(n830) );
  INV0 U552 ( .A(n176), .Q(n771) );
  INV0 U553 ( .A(n244), .Q(n819) );
  NOR22 U554 ( .A(A[7]), .B(B[7]), .Q(n252) );
  NOR22 U555 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NAND21 U556 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U557 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND20 U558 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND21 U559 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U560 ( .A(n39), .Q(n801) );
  NAND21 U561 ( .A(n793), .B(n62), .Q(n9) );
  NAND20 U562 ( .A(n829), .B(n275), .Q(n36) );
  XNR20 U563 ( .A(n34), .B(n828), .Q(SUM[4]) );
  NAND20 U564 ( .A(n830), .B(n272), .Q(n35) );
  INV3 U565 ( .A(n769), .Q(n777) );
  AOI211 U566 ( .A(n769), .B(n55), .C(n56), .Q(n54) );
  INV3 U567 ( .A(n219), .Q(n815) );
  INV0 U568 ( .A(n240), .Q(n818) );
  AOI211 U569 ( .A(n60), .B(n800), .C(n799), .Q(n47) );
  INV3 U570 ( .A(n51), .Q(n799) );
  NAND20 U571 ( .A(n171), .B(n779), .Q(n158) );
  INV3 U572 ( .A(n163), .Q(n780) );
  AOI210 U573 ( .A(n776), .B(n803), .C(n802), .Q(n141) );
  AOI210 U574 ( .A(n776), .B(n122), .C(n123), .Q(n121) );
  NAND22 U575 ( .A(n815), .B(n808), .Q(n208) );
  AOI210 U576 ( .A(n813), .B(n808), .C(n810), .Q(n209) );
  NOR21 U577 ( .A(n194), .B(n809), .Q(n190) );
  NAND20 U578 ( .A(n239), .B(n816), .Q(n226) );
  AOI210 U579 ( .A(n240), .B(n816), .C(n817), .Q(n227) );
  INV3 U580 ( .A(n231), .Q(n817) );
  NOR21 U581 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U582 ( .A(n788), .B(n792), .Q(n424) );
  INV3 U583 ( .A(n177), .Q(n778) );
  INV3 U584 ( .A(n212), .Q(n808) );
  INV3 U585 ( .A(n99), .Q(n792) );
  INV0 U586 ( .A(n70), .Q(n798) );
  INV0 U587 ( .A(n88), .Q(n796) );
  INV3 U588 ( .A(n126), .Q(n785) );
  INV3 U589 ( .A(n194), .Q(n807) );
  INV3 U590 ( .A(n107), .Q(n788) );
  INV3 U591 ( .A(n260), .Q(n825) );
  INV3 U592 ( .A(n61), .Q(n793) );
  INV3 U593 ( .A(n117), .Q(n784) );
  INV3 U594 ( .A(n241), .Q(n821) );
  INV3 U595 ( .A(n205), .Q(n812) );
  INV3 U596 ( .A(n137), .Q(n781) );
  INV3 U597 ( .A(n255), .Q(n823) );
  INV3 U598 ( .A(n252), .Q(n824) );
  INV3 U599 ( .A(n79), .Q(n797) );
  INV3 U600 ( .A(n185), .Q(n806) );
  NOR21 U601 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U602 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U603 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR22 U604 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR21 U605 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U606 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR21 U607 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND22 U608 ( .A(A[0]), .B(B[0]), .Q(n281) );
  INV3 U609 ( .A(n280), .Q(n834) );
  NOR21 U610 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U611 ( .A(n801), .B(n40), .Q(n7) );
  XNR21 U612 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U613 ( .A(n253), .B(n824), .Q(n31) );
  NAND20 U614 ( .A(n826), .B(n266), .Q(n34) );
  XNR21 U615 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NAND20 U616 ( .A(n798), .B(n71), .Q(n10) );
  NAND20 U617 ( .A(n792), .B(n100), .Q(n13) );
  XNR21 U618 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NAND20 U619 ( .A(n174), .B(n805), .Q(n21) );
  XNR21 U620 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U621 ( .A(n804), .B(n156), .Q(n19) );
  XNR21 U622 ( .A(n18), .B(n146), .Q(SUM[20]) );
  XNR21 U623 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND20 U624 ( .A(n785), .B(n127), .Q(n16) );
  XNR21 U625 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND20 U626 ( .A(n784), .B(n118), .Q(n15) );
  XNR21 U627 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NAND20 U628 ( .A(n796), .B(n89), .Q(n12) );
  XNR21 U629 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U630 ( .A(n812), .B(n206), .Q(n25) );
  XNR21 U631 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U632 ( .A(n807), .B(n195), .Q(n24) );
  NAND20 U633 ( .A(n771), .B(n177), .Q(n22) );
  XNR21 U634 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U635 ( .A(n816), .B(n231), .Q(n28) );
  XNR21 U636 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U637 ( .A(n224), .B(n814), .Q(n27) );
  NAND20 U638 ( .A(n819), .B(n245), .Q(n30) );
  XOR21 U639 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND20 U640 ( .A(n825), .B(n261), .Q(n33) );
  NAND20 U641 ( .A(n789), .B(n107), .Q(n14) );
  NAND20 U642 ( .A(n797), .B(n80), .Q(n11) );
  XNR21 U643 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND20 U644 ( .A(n779), .B(n163), .Q(n20) );
  XNR21 U645 ( .A(n17), .B(n139), .Q(SUM[21]) );
  NAND20 U646 ( .A(n781), .B(n138), .Q(n17) );
  XNR21 U647 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U648 ( .A(n806), .B(n186), .Q(n23) );
  XNR21 U649 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U650 ( .A(n821), .B(n242), .Q(n29) );
  XNR21 U651 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U652 ( .A(n808), .B(n213), .Q(n26) );
  XOR21 U653 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND20 U654 ( .A(n823), .B(n256), .Q(n32) );
  XNR21 U655 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XOR21 U656 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U657 ( .A(n831), .B(n279), .Q(n37) );
  XOR21 U658 ( .A(n36), .B(n832), .Q(SUM[2]) );
  INV3 U659 ( .A(n38), .Q(SUM[0]) );
  NAND22 U660 ( .A(n834), .B(n281), .Q(n38) );
endmodule


module adder_24 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_24_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module reg_7 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n5, n7, n9, n11, n13, n15, n17, n21, n23, n25, n27, n34, n49, n51,
         n53, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n55, n56, n57, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n103, n24, n26, n28, n29, n30, n32, n33,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n50, n52, n54, n101, n102, n104, n105, n106, n107, n108, n109, n110,
         n111, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328;

  DF3 Dout_reg_15_ ( .D(n74), .C(Clk), .Q(Dout[15]), .QN(n7) );
  DF3 Dout_reg_14_ ( .D(n75), .C(Clk), .Q(Dout[14]), .QN(n5) );
  DF3 Dout_reg_13_ ( .D(n87), .C(Clk), .Q(Dout[13]), .QN(n78) );
  DF3 Dout_reg_12_ ( .D(n88), .C(Clk), .Q(Dout[12]), .QN(n77) );
  DF3 Dout_reg_11_ ( .D(n89), .C(Clk), .Q(Dout[11]), .QN(n76) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n57) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n56) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n55) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n82) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n81) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n80) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n79) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n84) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n83) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n86) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n85) );
  DF3 Dout_reg_16_ ( .D(n73), .C(Clk), .Q(Dout[16]), .QN(n9) );
  DF3 Dout_reg_17_ ( .D(n72), .C(Clk), .Q(Dout[17]), .QN(n11) );
  DF3 Dout_reg_26_ ( .D(n63), .C(Clk), .Q(Dout[26]), .QN(n103) );
  DF3 Dout_reg_21_ ( .D(n68), .C(Clk), .Q(Dout[21]) );
  DF3 Dout_reg_18_ ( .D(n71), .C(Clk), .Q(Dout[18]), .QN(n13) );
  DF3 Dout_reg_25_ ( .D(n64), .C(Clk), .Q(Dout[25]), .QN(n27) );
  DF3 Dout_reg_22_ ( .D(n67), .C(Clk), .Q(Dout[22]), .QN(n21) );
  DF3 Dout_reg_24_ ( .D(n65), .C(Clk), .Q(Dout[24]), .QN(n25) );
  DF3 Dout_reg_23_ ( .D(n66), .C(Clk), .Q(Dout[23]), .QN(n23) );
  DF3 Dout_reg_19_ ( .D(n70), .C(Clk), .Q(Dout[19]), .QN(n15) );
  DF3 Dout_reg_20_ ( .D(n69), .C(Clk), .Q(Dout[20]), .QN(n17) );
  OAI212 U3 ( .A(n86), .B(n324), .C(n24), .Q(n99) );
  OAI212 U5 ( .A(n83), .B(n324), .C(n28), .Q(n98) );
  OAI212 U7 ( .A(n84), .B(n324), .C(n29), .Q(n97) );
  OAI212 U9 ( .A(n79), .B(n324), .C(n30), .Q(n96) );
  OAI212 U11 ( .A(n80), .B(n324), .C(n32), .Q(n95) );
  OAI212 U13 ( .A(n81), .B(n324), .C(n33), .Q(n94) );
  OAI212 U15 ( .A(n82), .B(n324), .C(n35), .Q(n93) );
  OAI212 U17 ( .A(n55), .B(n324), .C(n36), .Q(n92) );
  OAI212 U19 ( .A(n56), .B(n324), .C(n37), .Q(n91) );
  OAI212 U21 ( .A(n57), .B(n324), .C(n38), .Q(n90) );
  OAI212 U23 ( .A(n76), .B(n324), .C(n39), .Q(n89) );
  OAI212 U25 ( .A(n77), .B(n324), .C(n40), .Q(n88) );
  OAI212 U27 ( .A(n78), .B(n324), .C(n41), .Q(n87) );
  OAI212 U29 ( .A(n5), .B(n324), .C(n42), .Q(n75) );
  OAI212 U31 ( .A(n7), .B(n324), .C(n43), .Q(n74) );
  OAI212 U33 ( .A(n9), .B(n324), .C(n44), .Q(n73) );
  OAI212 U35 ( .A(n11), .B(n324), .C(n45), .Q(n72) );
  OAI212 U37 ( .A(n13), .B(n324), .C(n46), .Q(n71) );
  OAI212 U39 ( .A(n15), .B(n324), .C(n47), .Q(n70) );
  OAI212 U41 ( .A(n17), .B(n324), .C(n48), .Q(n69) );
  OAI212 U45 ( .A(n21), .B(n324), .C(n52), .Q(n67) );
  OAI212 U47 ( .A(n23), .B(n324), .C(n54), .Q(n66) );
  OAI212 U49 ( .A(n25), .B(n324), .C(n101), .Q(n65) );
  OAI212 U51 ( .A(n27), .B(n324), .C(n102), .Q(n64) );
  OAI212 U53 ( .A(n103), .B(n324), .C(n104), .Q(n63) );
  OAI212 U57 ( .A(n34), .B(n324), .C(n106), .Q(n61) );
  OAI212 U59 ( .A(n49), .B(n324), .C(n107), .Q(n60) );
  OAI212 U61 ( .A(n51), .B(n324), .C(n108), .Q(n59) );
  OAI212 U63 ( .A(n53), .B(n324), .C(n109), .Q(n58) );
  OAI212 U65 ( .A(n85), .B(n324), .C(n110), .Q(n100) );
  DF1 Dout_reg_31_ ( .D(n58), .C(Clk), .Q(Dout[31]), .QN(n53) );
  DF1 Dout_reg_30_ ( .D(n59), .C(Clk), .Q(Dout[30]), .QN(n51) );
  DF3 Dout_reg_29_ ( .D(n60), .C(Clk), .Q(Dout[29]), .QN(n49) );
  DF3 Dout_reg_28_ ( .D(n61), .C(Clk), .Q(Dout[28]), .QN(n34) );
  DF3 Dout_reg_27_ ( .D(n62), .C(Clk), .Q(Dout[27]) );
  NAND23 U4 ( .A(Din[28]), .B(n319), .Q(n106) );
  NAND23 U6 ( .A(Din[25]), .B(n320), .Q(n102) );
  NAND22 U8 ( .A(Dout[27]), .B(n111), .Q(n316) );
  NAND22 U10 ( .A(n105), .B(n316), .Q(n62) );
  NAND22 U12 ( .A(Dout[21]), .B(n111), .Q(n317) );
  NAND22 U14 ( .A(n317), .B(n50), .Q(n68) );
  NAND23 U16 ( .A(Din[21]), .B(n318), .Q(n50) );
  NAND23 U18 ( .A(Din[26]), .B(n319), .Q(n104) );
  NAND23 U20 ( .A(Din[29]), .B(n320), .Q(n107) );
  NAND23 U22 ( .A(Din[30]), .B(n319), .Q(n108) );
  NAND23 U24 ( .A(Din[31]), .B(n320), .Q(n109) );
  NAND23 U26 ( .A(Din[27]), .B(n320), .Q(n105) );
  CLKBU2 U28 ( .A(n325), .Q(n318) );
  CLKBU2 U30 ( .A(n326), .Q(n321) );
  CLKBU2 U32 ( .A(n326), .Q(n322) );
  CLKBU2 U34 ( .A(n326), .Q(n323) );
  CLKBU2 U36 ( .A(n325), .Q(n320) );
  CLKBU2 U38 ( .A(n325), .Q(n319) );
  CLKBU2 U40 ( .A(n26), .Q(n327) );
  INV3 U42 ( .A(n111), .Q(n324) );
  CLKBU2 U43 ( .A(n26), .Q(n325) );
  CLKBU2 U44 ( .A(n26), .Q(n326) );
  NAND22 U46 ( .A(Din[6]), .B(n327), .Q(n33) );
  NAND22 U48 ( .A(Din[7]), .B(n327), .Q(n35) );
  NAND22 U50 ( .A(Din[16]), .B(n322), .Q(n44) );
  NAND22 U52 ( .A(Din[17]), .B(n323), .Q(n45) );
  NAND22 U54 ( .A(Din[24]), .B(n318), .Q(n101) );
  NAND22 U55 ( .A(Din[20]), .B(n322), .Q(n48) );
  NAND22 U56 ( .A(Din[19]), .B(n323), .Q(n47) );
  NAND22 U58 ( .A(Din[18]), .B(n322), .Q(n46) );
  NAND22 U60 ( .A(Din[23]), .B(n318), .Q(n54) );
  NAND22 U62 ( .A(Din[22]), .B(n318), .Q(n52) );
  NAND22 U64 ( .A(Din[9]), .B(n321), .Q(n37) );
  NAND22 U66 ( .A(Din[10]), .B(n321), .Q(n38) );
  NAND22 U67 ( .A(Din[11]), .B(n321), .Q(n39) );
  NAND22 U68 ( .A(Din[12]), .B(n321), .Q(n40) );
  NAND22 U69 ( .A(Din[13]), .B(n323), .Q(n41) );
  NAND22 U70 ( .A(Din[14]), .B(n322), .Q(n42) );
  NAND22 U71 ( .A(Din[15]), .B(n323), .Q(n43) );
  NAND22 U72 ( .A(Din[8]), .B(n327), .Q(n36) );
  NAND22 U73 ( .A(Din[5]), .B(n327), .Q(n32) );
  NAND22 U74 ( .A(Din[2]), .B(n327), .Q(n28) );
  NAND22 U75 ( .A(Din[4]), .B(n327), .Q(n30) );
  NAND22 U76 ( .A(Din[3]), .B(n327), .Q(n29) );
  NOR21 U77 ( .A(n328), .B(Reset), .Q(n26) );
  INV3 U78 ( .A(Load), .Q(n328) );
  NAND22 U79 ( .A(Din[0]), .B(n319), .Q(n110) );
  NAND22 U80 ( .A(Din[1]), .B(n327), .Q(n24) );
  NOR20 U81 ( .A(Load), .B(Reset), .Q(n111) );
endmodule


module reg_6 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32,
         n35, n47, n49, n51, n53, n55, n57, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n58, n59, n60, n61, n62, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n103, n104, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396;

  DF3 Dout_reg_16_ ( .D(n78), .C(Clk), .Q(Dout[16]), .QN(n16) );
  DF3 Dout_reg_15_ ( .D(n79), .C(Clk), .Q(Dout[15]), .QN(n14) );
  DF3 Dout_reg_14_ ( .D(n80), .C(Clk), .Q(Dout[14]), .QN(n12) );
  DF3 Dout_reg_13_ ( .D(n81), .C(Clk), .Q(Dout[13]), .QN(n10) );
  DF3 Dout_reg_12_ ( .D(n82), .C(Clk), .Q(Dout[12]), .QN(n8) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n58) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n60) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n86) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n85) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n84) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n62) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n61) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n87) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n89) );
  DF3 Dout_reg_11_ ( .D(n83), .C(Clk), .Q(Dout[11]), .QN(n6) );
  DF3 Dout_reg_25_ ( .D(n69), .C(Clk), .Q(Dout[25]), .QN(n35) );
  DF3 Dout_reg_19_ ( .D(n75), .C(Clk), .Q(Dout[19]), .QN(n22) );
  DF3 Dout_reg_18_ ( .D(n76), .C(Clk), .Q(Dout[18]), .QN(n20) );
  DF3 Dout_reg_21_ ( .D(n73), .C(Clk), .Q(Dout[21]), .QN(n26) );
  DF3 Dout_reg_24_ ( .D(n70), .C(Clk), .Q(Dout[24]), .QN(n32) );
  DF3 Dout_reg_20_ ( .D(n74), .C(Clk), .Q(Dout[20]), .QN(n24) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n59) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n88) );
  DF3 Dout_reg_23_ ( .D(n71), .C(Clk), .Q(Dout[23]), .QN(n30) );
  DF3 Dout_reg_22_ ( .D(n72), .C(Clk), .Q(Dout[22]), .QN(n28) );
  DF3 Dout_reg_17_ ( .D(n77), .C(Clk), .Q(Dout[17]), .QN(n18) );
  OAI222 U3 ( .A(n88), .B(n361), .C(n363), .D(n395), .Q(n99) );
  OAI222 U4 ( .A(n87), .B(n361), .C(n362), .D(n394), .Q(n98) );
  OAI222 U5 ( .A(n61), .B(n361), .C(n103), .D(n393), .Q(n97) );
  OAI222 U6 ( .A(n62), .B(n361), .C(n363), .D(n390), .Q(n96) );
  OAI222 U7 ( .A(n84), .B(n361), .C(n362), .D(n391), .Q(n95) );
  OAI222 U8 ( .A(n85), .B(n361), .C(n103), .D(n392), .Q(n94) );
  OAI222 U9 ( .A(n86), .B(n361), .C(n363), .D(n389), .Q(n93) );
  OAI222 U10 ( .A(n60), .B(n361), .C(n362), .D(n387), .Q(n92) );
  OAI222 U11 ( .A(n59), .B(n361), .C(n103), .D(n388), .Q(n91) );
  OAI222 U12 ( .A(n58), .B(n361), .C(n363), .D(n386), .Q(n90) );
  OAI222 U13 ( .A(n6), .B(n361), .C(n362), .D(n379), .Q(n83) );
  OAI222 U14 ( .A(n8), .B(n361), .C(n103), .D(n383), .Q(n82) );
  OAI222 U15 ( .A(n10), .B(n361), .C(n363), .D(n381), .Q(n81) );
  OAI222 U16 ( .A(n12), .B(n361), .C(n362), .D(n382), .Q(n80) );
  OAI222 U17 ( .A(n14), .B(n361), .C(n103), .D(n380), .Q(n79) );
  OAI222 U18 ( .A(n16), .B(n361), .C(n363), .D(n384), .Q(n78) );
  OAI222 U19 ( .A(n18), .B(n361), .C(n362), .D(n385), .Q(n77) );
  OAI222 U20 ( .A(n20), .B(n361), .C(n103), .D(n378), .Q(n76) );
  OAI222 U21 ( .A(n22), .B(n361), .C(n363), .D(n377), .Q(n75) );
  OAI222 U22 ( .A(n24), .B(n361), .C(n362), .D(n376), .Q(n74) );
  OAI222 U23 ( .A(n26), .B(n361), .C(n103), .D(n374), .Q(n73) );
  OAI222 U24 ( .A(n28), .B(n361), .C(n375), .D(n363), .Q(n72) );
  OAI222 U25 ( .A(n30), .B(n361), .C(n362), .D(n371), .Q(n71) );
  OAI222 U26 ( .A(n32), .B(n361), .C(n103), .D(n372), .Q(n70) );
  OAI222 U27 ( .A(n35), .B(n361), .C(n363), .D(n373), .Q(n69) );
  OAI222 U28 ( .A(n47), .B(n361), .C(n362), .D(n370), .Q(n68) );
  OAI222 U29 ( .A(n49), .B(n361), .C(n103), .D(n369), .Q(n67) );
  OAI222 U30 ( .A(n51), .B(n361), .C(n363), .D(n368), .Q(n66) );
  OAI222 U31 ( .A(n53), .B(n361), .C(n362), .D(n367), .Q(n65) );
  OAI222 U32 ( .A(n55), .B(n361), .C(n103), .D(n366), .Q(n64) );
  OAI222 U33 ( .A(n57), .B(n361), .C(n363), .D(n365), .Q(n63) );
  OAI222 U34 ( .A(n89), .B(n361), .C(n362), .D(n396), .Q(n100) );
  DF1 Dout_reg_30_ ( .D(n64), .C(Clk), .Q(Dout[30]), .QN(n55) );
  DF1 Dout_reg_31_ ( .D(n63), .C(Clk), .Q(Dout[31]), .QN(n57) );
  DF1 Dout_reg_29_ ( .D(n65), .C(Clk), .Q(Dout[29]), .QN(n53) );
  DF3 Dout_reg_28_ ( .D(n66), .C(Clk), .Q(Dout[28]), .QN(n51) );
  DF1 Dout_reg_27_ ( .D(n67), .C(Clk), .Q(Dout[27]), .QN(n49) );
  DF1 Dout_reg_26_ ( .D(n68), .C(Clk), .Q(Dout[26]), .QN(n47) );
  INV3 U35 ( .A(Din[30]), .Q(n366) );
  INV3 U36 ( .A(Din[25]), .Q(n373) );
  INV3 U37 ( .A(Din[27]), .Q(n369) );
  INV2 U38 ( .A(Din[26]), .Q(n370) );
  INV3 U39 ( .A(Din[29]), .Q(n367) );
  INV3 U40 ( .A(Din[22]), .Q(n375) );
  INV3 U41 ( .A(Din[31]), .Q(n365) );
  INV3 U42 ( .A(Din[10]), .Q(n386) );
  INV3 U43 ( .A(Din[11]), .Q(n379) );
  INV3 U44 ( .A(Din[9]), .Q(n388) );
  INV3 U45 ( .A(Din[20]), .Q(n376) );
  INV3 U46 ( .A(Din[21]), .Q(n374) );
  INV6 U47 ( .A(Din[28]), .Q(n368) );
  CLKIN2 U48 ( .A(Din[8]), .Q(n387) );
  INV3 U49 ( .A(Din[23]), .Q(n371) );
  INV2 U50 ( .A(Din[7]), .Q(n389) );
  INV3 U51 ( .A(Din[17]), .Q(n385) );
  CLKIN3 U52 ( .A(Din[18]), .Q(n378) );
  INV2 U53 ( .A(Din[19]), .Q(n377) );
  INV2 U54 ( .A(Din[16]), .Q(n384) );
  INV2 U55 ( .A(Din[24]), .Q(n372) );
  INV2 U56 ( .A(Din[13]), .Q(n381) );
  INV2 U57 ( .A(Din[14]), .Q(n382) );
  CLKIN3 U58 ( .A(Din[5]), .Q(n391) );
  CLKIN2 U59 ( .A(Din[4]), .Q(n390) );
  INV2 U60 ( .A(Din[15]), .Q(n380) );
  INV2 U61 ( .A(Din[12]), .Q(n383) );
  CLKIN2 U62 ( .A(Din[6]), .Q(n392) );
  NAND22 U63 ( .A(n364), .B(n361), .Q(n362) );
  NAND22 U64 ( .A(n364), .B(n361), .Q(n363) );
  NAND22 U65 ( .A(n364), .B(n361), .Q(n103) );
  INV3 U66 ( .A(Reset), .Q(n364) );
  INV3 U67 ( .A(n104), .Q(n361) );
  INV3 U68 ( .A(Din[1]), .Q(n395) );
  INV3 U69 ( .A(Din[3]), .Q(n393) );
  INV3 U70 ( .A(Din[2]), .Q(n394) );
  INV3 U71 ( .A(Din[0]), .Q(n396) );
  NOR21 U72 ( .A(Load), .B(Reset), .Q(n104) );
endmodule


module adder_23_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n416, n490,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U77 ( .A(n91), .B(n754), .C(n92), .Q(n90) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n754), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n758), .B(n754), .C(n755), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U189 ( .A(n176), .B(n754), .C(n177), .Q(n175) );
  AOI212 U195 ( .A(n490), .B(n179), .C(n180), .Q(n178) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n268), .B(n248), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U448 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U418 ( .A(n102), .B(n754), .C(n103), .Q(n101) );
  OAI212 U421 ( .A(n129), .B(n754), .C(n130), .Q(n128) );
  OAI212 U435 ( .A(n140), .B(n754), .C(n141), .Q(n139) );
  OAI212 U427 ( .A(n82), .B(n754), .C(n83), .Q(n81) );
  OAI212 U609 ( .A(n760), .B(n754), .C(n753), .Q(n108) );
  OAI212 U611 ( .A(n73), .B(n754), .C(n74), .Q(n72) );
  OAI212 U353 ( .A(n226), .B(n776), .C(n227), .Q(n225) );
  OAI212 U385 ( .A(n208), .B(n776), .C(n209), .Q(n207) );
  OAI212 U414 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  AOI212 U415 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U387 ( .A(n774), .B(n776), .C(n772), .Q(n232) );
  OAI212 U395 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U401 ( .A(n194), .B(n763), .C(n195), .Q(n191) );
  OAI212 U405 ( .A(n244), .B(n776), .C(n245), .Q(n243) );
  OAI212 U429 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U439 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U457 ( .A(n197), .B(n776), .C(n198), .Q(n196) );
  OAI212 U428 ( .A(n42), .B(n754), .C(n43), .Q(n41) );
  OAI212 U430 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U360 ( .A(n53), .B(n754), .C(n54), .Q(n52) );
  OAI212 U497 ( .A(n813), .B(n5), .C(n814), .Q(n56) );
  OAI212 U451 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  AOI212 U423 ( .A(n240), .B(n221), .C(n222), .Q(n416) );
  OAI212 U436 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI212 U478 ( .A(n88), .B(n788), .C(n89), .Q(n85) );
  OAI212 U488 ( .A(n151), .B(n754), .C(n152), .Q(n146) );
  NAND22 U349 ( .A(n771), .B(n203), .Q(n197) );
  NAND22 U350 ( .A(A[24]), .B(B[24]), .Q(n107) );
  XNR22 U351 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND22 U352 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND22 U354 ( .A(n111), .B(n66), .Q(n64) );
  CLKIN6 U355 ( .A(n112), .Q(n751) );
  INV12 U356 ( .A(n751), .Q(n752) );
  NOR22 U357 ( .A(B[12]), .B(A[12]), .Q(n212) );
  AOI212 U358 ( .A(n752), .B(n84), .C(n85), .Q(n83) );
  AOI212 U359 ( .A(n752), .B(n97), .C(n98), .Q(n92) );
  INV1 U361 ( .A(n752), .Q(n753) );
  NOR23 U362 ( .A(n79), .B(n88), .Q(n77) );
  NOR24 U363 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND21 U364 ( .A(A[27]), .B(B[27]), .Q(n80) );
  XNR22 U365 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND26 U366 ( .A(n258), .B(n250), .Q(n248) );
  NOR24 U367 ( .A(n252), .B(n255), .Q(n250) );
  NOR22 U368 ( .A(n173), .B(n176), .Q(n171) );
  NOR22 U369 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR23 U370 ( .A(n99), .B(n106), .Q(n97) );
  NOR22 U371 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR23 U372 ( .A(n205), .B(n212), .Q(n203) );
  NOR22 U373 ( .A(n271), .B(n274), .Q(n269) );
  NAND22 U374 ( .A(n97), .B(n77), .Q(n6) );
  NAND22 U375 ( .A(n135), .B(n115), .Q(n113) );
  NOR22 U376 ( .A(n155), .B(n162), .Q(n153) );
  AOI211 U377 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR22 U378 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND22 U379 ( .A(n759), .B(n801), .Q(n140) );
  NAND22 U380 ( .A(n171), .B(n153), .Q(n151) );
  NOR23 U381 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NOR22 U382 ( .A(B[15]), .B(A[15]), .Q(n185) );
  XNR21 U383 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR21 U384 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR21 U386 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR21 U388 ( .A(n12), .B(n90), .Q(SUM[26]) );
  AOI211 U389 ( .A(n781), .B(n779), .C(n780), .Q(n262) );
  XOR21 U390 ( .A(n32), .B(n257), .Q(SUM[6]) );
  XNR21 U391 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XNR21 U392 ( .A(n26), .B(n214), .Q(SUM[12]) );
  XNR21 U393 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND21 U394 ( .A(n803), .B(n242), .Q(n29) );
  NAND21 U396 ( .A(n761), .B(n186), .Q(n23) );
  NAND23 U397 ( .A(n203), .B(n183), .Q(n181) );
  NOR22 U398 ( .A(B[1]), .B(A[1]), .Q(n278) );
  XOR22 U399 ( .A(n22), .B(n754), .Q(SUM[16]) );
  NOR22 U400 ( .A(n260), .B(n265), .Q(n258) );
  NOR24 U402 ( .A(n223), .B(n230), .Q(n221) );
  AOI212 U403 ( .A(n781), .B(n258), .C(n259), .Q(n257) );
  INV3 U404 ( .A(n268), .Q(n781) );
  NAND22 U406 ( .A(A[17]), .B(B[17]), .Q(n174) );
  XNR22 U407 ( .A(n225), .B(n27), .Q(SUM[11]) );
  XNR22 U408 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NOR23 U409 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NOR24 U410 ( .A(B[14]), .B(A[14]), .Q(n194) );
  XNR22 U411 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NAND22 U412 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U413 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NOR23 U416 ( .A(B[3]), .B(A[3]), .Q(n271) );
  XNR22 U417 ( .A(n19), .B(n157), .Q(SUM[19]) );
  XNR22 U419 ( .A(n23), .B(n187), .Q(SUM[15]) );
  INV10 U420 ( .A(n247), .Q(n776) );
  OAI212 U422 ( .A(n219), .B(n776), .C(n416), .Q(n214) );
  OAI211 U424 ( .A(n188), .B(n776), .C(n189), .Q(n187) );
  OAI212 U425 ( .A(n268), .B(n248), .C(n249), .Q(n490) );
  XNR22 U426 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XNR22 U431 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND22 U432 ( .A(A[16]), .B(B[16]), .Q(n177) );
  XNR22 U433 ( .A(n21), .B(n175), .Q(SUM[17]) );
  AOI212 U434 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NAND24 U437 ( .A(n239), .B(n221), .Q(n219) );
  NOR22 U438 ( .A(n241), .B(n244), .Q(n239) );
  INV6 U440 ( .A(n219), .Q(n771) );
  XOR20 U441 ( .A(n36), .B(n785), .Q(SUM[2]) );
  OAI211 U442 ( .A(n274), .B(n785), .C(n275), .Q(n273) );
  INV3 U443 ( .A(n277), .Q(n785) );
  NOR22 U444 ( .A(n185), .B(n194), .Q(n183) );
  XNR22 U445 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U446 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND21 U447 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND22 U449 ( .A(n111), .B(n97), .Q(n91) );
  NOR24 U450 ( .A(n113), .B(n151), .Q(n111) );
  OAI212 U452 ( .A(n120), .B(n754), .C(n121), .Q(n119) );
  NOR23 U453 ( .A(B[10]), .B(A[10]), .Q(n230) );
  OAI212 U454 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  NOR23 U455 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND21 U456 ( .A(n806), .B(n127), .Q(n16) );
  OAI211 U458 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI211 U459 ( .A(n126), .B(n798), .C(n127), .Q(n123) );
  NAND21 U460 ( .A(A[22]), .B(B[22]), .Q(n127) );
  BUF15 U461 ( .A(n178), .Q(n754) );
  INV2 U462 ( .A(n135), .Q(n797) );
  NAND22 U463 ( .A(n759), .B(n135), .Q(n129) );
  NOR22 U464 ( .A(n137), .B(n144), .Q(n135) );
  NAND22 U465 ( .A(n759), .B(n122), .Q(n120) );
  AOI211 U466 ( .A(n756), .B(n122), .C(n123), .Q(n121) );
  NOR21 U467 ( .A(n126), .B(n797), .Q(n122) );
  CLKIN3 U468 ( .A(n145), .Q(n802) );
  INV4 U469 ( .A(n151), .Q(n759) );
  NAND21 U470 ( .A(n111), .B(n792), .Q(n73) );
  NAND21 U471 ( .A(n55), .B(n111), .Q(n53) );
  NAND21 U472 ( .A(n111), .B(n44), .Q(n42) );
  NAND22 U473 ( .A(n111), .B(n84), .Q(n82) );
  CLKIN2 U474 ( .A(n111), .Q(n760) );
  OAI211 U475 ( .A(n64), .B(n754), .C(n65), .Q(n63) );
  XNR22 U476 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND21 U477 ( .A(n111), .B(n800), .Q(n102) );
  INV0 U479 ( .A(n106), .Q(n800) );
  CLKIN1 U480 ( .A(n136), .Q(n798) );
  INV0 U481 ( .A(n204), .Q(n763) );
  AOI211 U482 ( .A(n769), .B(n190), .C(n191), .Q(n189) );
  NAND21 U483 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND20 U484 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND21 U485 ( .A(A[9]), .B(B[9]), .Q(n242) );
  AOI211 U486 ( .A(n752), .B(n66), .C(n67), .Q(n65) );
  INV0 U487 ( .A(n255), .Q(n777) );
  NAND20 U489 ( .A(n812), .B(n62), .Q(n9) );
  NAND20 U490 ( .A(n800), .B(n107), .Q(n14) );
  AOI211 U491 ( .A(n221), .B(n240), .C(n222), .Q(n220) );
  NAND20 U492 ( .A(n808), .B(n89), .Q(n12) );
  NAND20 U493 ( .A(n809), .B(n174), .Q(n21) );
  AOI211 U494 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  XOR21 U495 ( .A(n30), .B(n776), .Q(SUM[8]) );
  NAND20 U496 ( .A(n816), .B(n71), .Q(n10) );
  NAND20 U498 ( .A(n790), .B(n100), .Q(n13) );
  NAND20 U499 ( .A(n805), .B(n118), .Q(n15) );
  INV0 U500 ( .A(n274), .Q(n783) );
  INV0 U501 ( .A(n271), .Q(n782) );
  INV0 U502 ( .A(n252), .Q(n775) );
  INV0 U503 ( .A(n194), .Q(n762) );
  INV0 U504 ( .A(n278), .Q(n804) );
  NAND21 U505 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND21 U506 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NAND22 U507 ( .A(A[8]), .B(B[8]), .Q(n245) );
  INV3 U508 ( .A(n416), .Q(n769) );
  NOR20 U509 ( .A(n813), .B(n6), .Q(n55) );
  INV0 U510 ( .A(n6), .Q(n792) );
  INV3 U511 ( .A(n152), .Q(n756) );
  AOI210 U512 ( .A(n769), .B(n203), .C(n204), .Q(n198) );
  AOI210 U513 ( .A(n756), .B(n135), .C(n136), .Q(n130) );
  NOR23 U514 ( .A(n181), .B(n219), .Q(n179) );
  NOR20 U515 ( .A(n46), .B(n6), .Q(n44) );
  NAND21 U516 ( .A(n771), .B(n190), .Q(n188) );
  NAND20 U517 ( .A(n171), .B(n795), .Q(n158) );
  NAND20 U518 ( .A(n239), .B(n770), .Q(n226) );
  CLKIN3 U519 ( .A(n59), .Q(n813) );
  INV0 U520 ( .A(n88), .Q(n808) );
  INV0 U521 ( .A(n176), .Q(n757) );
  INV0 U522 ( .A(n173), .Q(n809) );
  NAND20 U523 ( .A(n762), .B(n195), .Q(n24) );
  INV0 U524 ( .A(n213), .Q(n767) );
  INV0 U525 ( .A(n61), .Q(n812) );
  INV0 U526 ( .A(n99), .Q(n790) );
  NAND20 U527 ( .A(n801), .B(n145), .Q(n18) );
  INV0 U528 ( .A(n205), .Q(n764) );
  INV0 U529 ( .A(n185), .Q(n761) );
  INV0 U530 ( .A(n126), .Q(n806) );
  CLKIN0 U531 ( .A(n171), .Q(n758) );
  NAND20 U532 ( .A(n795), .B(n163), .Q(n20) );
  INV0 U533 ( .A(n117), .Q(n805) );
  NAND20 U534 ( .A(n777), .B(n256), .Q(n32) );
  INV0 U535 ( .A(n231), .Q(n768) );
  CLKIN0 U536 ( .A(n203), .Q(n765) );
  XOR20 U537 ( .A(n281), .B(n37), .Q(SUM[1]) );
  INV0 U538 ( .A(n244), .Q(n773) );
  NAND20 U539 ( .A(n783), .B(n275), .Q(n36) );
  INV0 U540 ( .A(n260), .Q(n778) );
  CLKIN2 U541 ( .A(n97), .Q(n791) );
  XNR20 U542 ( .A(n34), .B(n781), .Q(SUM[4]) );
  NAND20 U543 ( .A(n779), .B(n266), .Q(n34) );
  INV0 U544 ( .A(n241), .Q(n803) );
  CLKIN0 U545 ( .A(n239), .Q(n774) );
  NAND20 U546 ( .A(n770), .B(n231), .Q(n28) );
  OAI210 U547 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND20 U548 ( .A(n782), .B(n272), .Q(n35) );
  NAND20 U549 ( .A(n59), .B(n810), .Q(n46) );
  NAND20 U550 ( .A(n775), .B(n253), .Q(n31) );
  INV0 U551 ( .A(n70), .Q(n816) );
  INV0 U552 ( .A(n223), .Q(n787) );
  NAND20 U553 ( .A(n766), .B(n213), .Q(n26) );
  INV0 U554 ( .A(n266), .Q(n780) );
  NAND21 U555 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NOR22 U556 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR22 U557 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR22 U558 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR22 U559 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U560 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR21 U561 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR21 U562 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NAND21 U563 ( .A(B[1]), .B(A[1]), .Q(n279) );
  NAND20 U564 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U565 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U566 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND21 U567 ( .A(A[25]), .B(B[25]), .Q(n100) );
  AOI210 U568 ( .A(n752), .B(n55), .C(n56), .Q(n54) );
  INV3 U569 ( .A(n60), .Q(n814) );
  AOI210 U570 ( .A(n752), .B(n792), .C(n789), .Q(n74) );
  CLKIN0 U571 ( .A(n5), .Q(n789) );
  INV0 U572 ( .A(n240), .Q(n772) );
  NAND22 U573 ( .A(n771), .B(n766), .Q(n208) );
  INV0 U574 ( .A(n172), .Q(n755) );
  NAND22 U575 ( .A(n807), .B(n80), .Q(n11) );
  INV3 U576 ( .A(n79), .Q(n807) );
  NAND22 U577 ( .A(n279), .B(n804), .Q(n37) );
  XOR21 U578 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND22 U579 ( .A(n778), .B(n261), .Q(n33) );
  NAND22 U580 ( .A(n757), .B(n177), .Q(n22) );
  NAND22 U581 ( .A(n773), .B(n245), .Q(n30) );
  NAND22 U582 ( .A(n787), .B(n224), .Q(n27) );
  XNR21 U583 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U584 ( .A(n793), .B(n156), .Q(n19) );
  INV3 U585 ( .A(n155), .Q(n793) );
  NAND22 U586 ( .A(n764), .B(n206), .Q(n25) );
  XNR21 U587 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR21 U588 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND22 U589 ( .A(n810), .B(n51), .Q(n8) );
  NAND22 U590 ( .A(n796), .B(n138), .Q(n17) );
  INV3 U591 ( .A(n137), .Q(n796) );
  NOR21 U592 ( .A(n61), .B(n70), .Q(n59) );
  NOR21 U593 ( .A(n70), .B(n6), .Q(n66) );
  NOR21 U594 ( .A(n117), .B(n126), .Q(n115) );
  AOI210 U595 ( .A(n240), .B(n770), .C(n768), .Q(n227) );
  AOI210 U596 ( .A(n172), .B(n795), .C(n794), .Q(n159) );
  INV3 U597 ( .A(n163), .Q(n794) );
  INV0 U598 ( .A(n98), .Q(n788) );
  AOI210 U599 ( .A(n752), .B(n44), .C(n45), .Q(n43) );
  AOI211 U600 ( .A(n60), .B(n810), .C(n811), .Q(n47) );
  INV3 U601 ( .A(n51), .Q(n811) );
  AOI211 U602 ( .A(n752), .B(n800), .C(n799), .Q(n103) );
  INV3 U603 ( .A(n107), .Q(n799) );
  AOI211 U604 ( .A(n769), .B(n766), .C(n767), .Q(n209) );
  AOI211 U605 ( .A(n756), .B(n801), .C(n802), .Q(n141) );
  INV3 U606 ( .A(n144), .Q(n801) );
  INV3 U607 ( .A(n162), .Q(n795) );
  INV3 U608 ( .A(n212), .Q(n766) );
  INV3 U610 ( .A(n230), .Q(n770) );
  NOR21 U612 ( .A(n88), .B(n791), .Q(n84) );
  NOR21 U613 ( .A(n194), .B(n765), .Q(n190) );
  INV3 U614 ( .A(n265), .Q(n779) );
  NOR21 U615 ( .A(B[28]), .B(A[28]), .Q(n70) );
  XNR21 U616 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U617 ( .A(n815), .B(n40), .Q(n7) );
  NAND22 U618 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR22 U619 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR21 U620 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR22 U621 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR22 U622 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR22 U623 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR22 U624 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR22 U625 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U626 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND22 U627 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND22 U628 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U629 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND22 U630 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND22 U631 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U632 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND22 U633 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND22 U634 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U635 ( .A(A[7]), .B(B[7]), .Q(n253) );
  INV3 U636 ( .A(n38), .Q(SUM[0]) );
  NAND20 U637 ( .A(n786), .B(n281), .Q(n38) );
  INV3 U638 ( .A(n280), .Q(n786) );
  NOR20 U639 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U640 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U641 ( .A(n50), .Q(n810) );
  NOR21 U642 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U643 ( .A(n39), .Q(n815) );
  NOR21 U644 ( .A(B[31]), .B(A[31]), .Q(n39) );
endmodule


module adder_23 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_23_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_22_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n419, n420, n421,
         n426, n432, n500, n504, n508, n575, n593, n596, n666, n678, n680,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n825, n826, n827;

  OAI212 U11 ( .A(n42), .B(n758), .C(n43), .Q(n41) );
  OAI212 U135 ( .A(n137), .B(n145), .C(n138), .Q(n136) );
  AOI212 U157 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n825), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U416 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U483 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  AOI212 U537 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI212 U448 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U412 ( .A(n821), .B(n813), .C(n819), .Q(n232) );
  OAI212 U413 ( .A(n226), .B(n813), .C(n227), .Q(n225) );
  OAI212 U414 ( .A(n197), .B(n813), .C(n198), .Q(n196) );
  OAI212 U505 ( .A(n194), .B(n807), .C(n195), .Q(n191) );
  NOR24 U364 ( .A(B[26]), .B(A[26]), .Q(n88) );
  OAI212 U418 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  OAI212 U517 ( .A(n91), .B(n758), .C(n92), .Q(n90) );
  NOR24 U536 ( .A(n79), .B(n88), .Q(n77) );
  OAI212 U544 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U550 ( .A(n152), .B(n113), .C(n114), .Q(n112) );
  OAI212 U556 ( .A(n88), .B(n776), .C(n89), .Q(n85) );
  NOR23 U349 ( .A(n144), .B(n137), .Q(n135) );
  NOR23 U350 ( .A(B[21]), .B(A[21]), .Q(n137) );
  CLKIN6 U351 ( .A(n155), .Q(n756) );
  XNR22 U352 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U353 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND24 U354 ( .A(n153), .B(n171), .Q(n151) );
  NAND26 U355 ( .A(n203), .B(n183), .Q(n181) );
  NOR24 U356 ( .A(n185), .B(n194), .Q(n183) );
  NOR24 U357 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR24 U358 ( .A(B[18]), .B(A[18]), .Q(n162) );
  AOI212 U359 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  AOI211 U360 ( .A(n60), .B(n760), .C(n761), .Q(n47) );
  NAND24 U361 ( .A(n500), .B(n103), .Q(n101) );
  NAND28 U362 ( .A(n115), .B(n135), .Q(n113) );
  NOR23 U363 ( .A(A[20]), .B(B[20]), .Q(n144) );
  INV3 U365 ( .A(n84), .Q(n779) );
  NOR22 U366 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR23 U367 ( .A(A[11]), .B(B[11]), .Q(n223) );
  INV3 U368 ( .A(n106), .Q(n778) );
  NAND23 U369 ( .A(n752), .B(n756), .Q(n757) );
  NOR23 U370 ( .A(n223), .B(n230), .Q(n221) );
  NOR22 U371 ( .A(A[29]), .B(B[29]), .Q(n61) );
  NAND23 U372 ( .A(n55), .B(n111), .Q(n53) );
  NOR23 U373 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NAND22 U374 ( .A(n111), .B(n778), .Q(n102) );
  NOR23 U375 ( .A(n173), .B(n176), .Q(n171) );
  INV3 U376 ( .A(n151), .Q(n790) );
  NAND26 U377 ( .A(n419), .B(n100), .Q(n98) );
  NOR21 U378 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR22 U379 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR22 U380 ( .A(A[10]), .B(B[10]), .Q(n230) );
  NOR23 U381 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NAND23 U382 ( .A(n775), .B(n797), .Q(n593) );
  NAND22 U383 ( .A(n768), .B(n80), .Q(n11) );
  NAND22 U384 ( .A(A[16]), .B(B[16]), .Q(n177) );
  AOI211 U385 ( .A(n812), .B(n258), .C(n259), .Q(n257) );
  NAND22 U386 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND22 U387 ( .A(B[10]), .B(A[10]), .Q(n231) );
  NAND22 U388 ( .A(B[12]), .B(A[12]), .Q(n213) );
  NAND22 U389 ( .A(B[14]), .B(A[14]), .Q(n195) );
  XNR21 U390 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR21 U391 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NOR23 U392 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NAND23 U393 ( .A(n757), .B(n156), .Q(n154) );
  CLKBU15 U394 ( .A(n178), .Q(n758) );
  INV1 U395 ( .A(n789), .Q(n751) );
  NOR24 U396 ( .A(A[17]), .B(B[17]), .Q(n173) );
  OAI212 U397 ( .A(n758), .B(n129), .C(n130), .Q(n128) );
  XNR22 U398 ( .A(n17), .B(n139), .Q(SUM[21]) );
  OAI212 U399 ( .A(n140), .B(n758), .C(n141), .Q(n139) );
  OAI212 U400 ( .A(n758), .B(n120), .C(n121), .Q(n119) );
  INV6 U401 ( .A(n163), .Q(n752) );
  CLKIN1 U402 ( .A(n752), .Q(n753) );
  AOI212 U403 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NAND22 U404 ( .A(A[6]), .B(B[6]), .Q(n256) );
  INV2 U405 ( .A(n152), .Q(n789) );
  NOR22 U406 ( .A(n88), .B(n780), .Q(n84) );
  NAND22 U407 ( .A(n790), .B(n122), .Q(n120) );
  NAND22 U408 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NOR23 U409 ( .A(B[14]), .B(A[14]), .Q(n194) );
  INV1 U410 ( .A(n220), .Q(n796) );
  OAI210 U411 ( .A(n219), .B(n813), .C(n220), .Q(n214) );
  AOI210 U415 ( .A(n796), .B(n203), .C(n420), .Q(n198) );
  NOR24 U417 ( .A(n181), .B(n219), .Q(n179) );
  OAI211 U419 ( .A(n89), .B(n79), .C(n80), .Q(n426) );
  NAND23 U420 ( .A(n763), .B(n797), .Q(n666) );
  INV3 U421 ( .A(n53), .Q(n763) );
  CLKIN2 U422 ( .A(n421), .Q(n767) );
  OAI211 U423 ( .A(n126), .B(n784), .C(n127), .Q(n123) );
  NOR23 U424 ( .A(B[30]), .B(A[30]), .Q(n50) );
  CLKIN3 U425 ( .A(n162), .Q(n792) );
  NAND22 U426 ( .A(B[17]), .B(A[17]), .Q(n174) );
  NAND26 U427 ( .A(n508), .B(n186), .Q(n184) );
  NAND24 U428 ( .A(n803), .B(n802), .Q(n508) );
  INV0 U429 ( .A(n205), .Q(n805) );
  NAND21 U430 ( .A(n781), .B(n89), .Q(n12) );
  OAI212 U431 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  CLKIN15 U432 ( .A(n754), .Q(n755) );
  NOR22 U433 ( .A(n244), .B(n241), .Q(n239) );
  XNR22 U434 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NAND23 U435 ( .A(n596), .B(n74), .Q(n72) );
  NAND20 U436 ( .A(n171), .B(n792), .Q(n158) );
  NAND21 U437 ( .A(B[11]), .B(A[11]), .Q(n224) );
  NAND21 U438 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND23 U439 ( .A(A[26]), .B(B[26]), .Q(n89) );
  OAI211 U440 ( .A(n158), .B(n758), .C(n159), .Q(n157) );
  OAI211 U441 ( .A(n794), .B(n758), .C(n795), .Q(n164) );
  INV1 U442 ( .A(n60), .Q(n765) );
  NAND21 U443 ( .A(B[19]), .B(A[19]), .Q(n156) );
  OAI211 U444 ( .A(n213), .B(n205), .C(n206), .Q(n420) );
  INV6 U445 ( .A(n755), .Q(n771) );
  NOR24 U446 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NAND26 U447 ( .A(n83), .B(n593), .Q(n81) );
  CLKIN6 U449 ( .A(n575), .Q(n782) );
  NAND22 U450 ( .A(n797), .B(n774), .Q(n500) );
  AOI212 U451 ( .A(n755), .B(n778), .C(n777), .Q(n103) );
  NOR24 U452 ( .A(n117), .B(n126), .Q(n115) );
  INV3 U453 ( .A(n102), .Q(n774) );
  AOI212 U454 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  CLKIN3 U455 ( .A(n247), .Q(n813) );
  INV0 U456 ( .A(n753), .Q(n791) );
  XNR22 U457 ( .A(n10), .B(n72), .Q(SUM[28]) );
  AOI210 U458 ( .A(n789), .B(n788), .C(n787), .Q(n141) );
  NAND20 U459 ( .A(n790), .B(n788), .Q(n140) );
  INV1 U460 ( .A(n144), .Q(n788) );
  NAND22 U461 ( .A(n111), .B(n66), .Q(n64) );
  AOI212 U462 ( .A(n755), .B(n97), .C(n98), .Q(n92) );
  OAI211 U463 ( .A(n208), .B(n813), .C(n209), .Q(n207) );
  OAI211 U464 ( .A(n188), .B(n813), .C(n189), .Q(n187) );
  NAND24 U465 ( .A(n59), .B(n760), .Q(n46) );
  INV6 U466 ( .A(n112), .Q(n754) );
  INV3 U467 ( .A(n135), .Q(n786) );
  XOR20 U468 ( .A(n32), .B(n257), .Q(SUM[6]) );
  AOI210 U469 ( .A(n812), .B(n814), .C(n815), .Q(n262) );
  OAI211 U470 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NAND21 U471 ( .A(A[3]), .B(B[3]), .Q(n272) );
  OAI212 U472 ( .A(n773), .B(n758), .C(n771), .Q(n108) );
  XNR22 U473 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NAND22 U474 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV3 U475 ( .A(n111), .Q(n773) );
  NAND22 U476 ( .A(n111), .B(n770), .Q(n73) );
  NAND22 U477 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND24 U478 ( .A(n666), .B(n54), .Q(n52) );
  AOI212 U479 ( .A(n98), .B(n77), .C(n78), .Q(n678) );
  NAND21 U480 ( .A(A[30]), .B(B[30]), .Q(n51) );
  OAI212 U481 ( .A(n5), .B(n46), .C(n47), .Q(n45) );
  NOR21 U482 ( .A(n126), .B(n786), .Q(n122) );
  NOR24 U484 ( .A(n46), .B(n6), .Q(n44) );
  AOI212 U485 ( .A(n755), .B(n770), .C(n767), .Q(n74) );
  CLKIN1 U486 ( .A(n241), .Q(n820) );
  NAND28 U487 ( .A(n97), .B(n77), .Q(n6) );
  CLKIN6 U488 ( .A(n97), .Q(n780) );
  NOR24 U489 ( .A(n575), .B(n106), .Q(n97) );
  NOR23 U490 ( .A(n70), .B(n6), .Q(n66) );
  NOR23 U491 ( .A(n764), .B(n6), .Q(n55) );
  INV6 U492 ( .A(n6), .Q(n770) );
  INV1 U493 ( .A(n61), .Q(n762) );
  INV0 U494 ( .A(n79), .Q(n768) );
  NAND21 U495 ( .A(n51), .B(n760), .Q(n8) );
  NOR24 U496 ( .A(n779), .B(n771), .Q(n680) );
  NOR24 U497 ( .A(n85), .B(n680), .Q(n83) );
  NAND24 U498 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NOR24 U499 ( .A(A[25]), .B(B[25]), .Q(n575) );
  XNR22 U500 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND24 U501 ( .A(n782), .B(n777), .Q(n419) );
  AOI212 U502 ( .A(n755), .B(n44), .C(n45), .Q(n43) );
  OAI211 U503 ( .A(n151), .B(n758), .C(n751), .Q(n146) );
  AOI212 U504 ( .A(n755), .B(n55), .C(n56), .Q(n54) );
  OAI212 U506 ( .A(n678), .B(n70), .C(n71), .Q(n67) );
  AOI212 U507 ( .A(n755), .B(n66), .C(n67), .Q(n65) );
  AOI212 U508 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR24 U509 ( .A(n252), .B(n255), .Q(n250) );
  NOR22 U510 ( .A(B[6]), .B(A[6]), .Q(n255) );
  XNR22 U511 ( .A(n11), .B(n81), .Q(SUM[27]) );
  INV3 U512 ( .A(n136), .Q(n784) );
  OAI211 U513 ( .A(n176), .B(n758), .C(n177), .Q(n175) );
  OAI212 U514 ( .A(n241), .B(n245), .C(n242), .Q(n240) );
  OAI210 U515 ( .A(n245), .B(n241), .C(n242), .Q(n504) );
  NAND22 U516 ( .A(B[9]), .B(A[9]), .Q(n242) );
  AOI210 U518 ( .A(n789), .B(n135), .C(n136), .Q(n130) );
  NAND21 U519 ( .A(B[23]), .B(A[23]), .Q(n118) );
  CLKIN4 U520 ( .A(n59), .Q(n764) );
  NOR22 U521 ( .A(n61), .B(n70), .Q(n59) );
  NAND26 U522 ( .A(n239), .B(n221), .Q(n219) );
  NAND21 U523 ( .A(n790), .B(n135), .Q(n129) );
  NOR23 U524 ( .A(B[28]), .B(A[28]), .Q(n70) );
  INV1 U525 ( .A(n98), .Q(n776) );
  NAND21 U526 ( .A(B[15]), .B(A[15]), .Q(n186) );
  INV10 U527 ( .A(n758), .Q(n797) );
  NAND21 U528 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND22 U529 ( .A(B[20]), .B(A[20]), .Q(n145) );
  NAND21 U530 ( .A(A[13]), .B(B[13]), .Q(n206) );
  XNR22 U531 ( .A(n9), .B(n63), .Q(SUM[29]) );
  OAI212 U532 ( .A(n64), .B(n758), .C(n65), .Q(n63) );
  NOR24 U533 ( .A(A[19]), .B(B[19]), .Q(n155) );
  OAI210 U534 ( .A(n244), .B(n813), .C(n245), .Q(n243) );
  AOI212 U535 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  NOR23 U538 ( .A(n162), .B(n155), .Q(n153) );
  XNR22 U539 ( .A(n7), .B(n41), .Q(SUM[31]) );
  INV2 U540 ( .A(n203), .Q(n806) );
  NAND22 U541 ( .A(n799), .B(n203), .Q(n197) );
  NOR24 U542 ( .A(n212), .B(n205), .Q(n203) );
  AOI212 U543 ( .A(n98), .B(n77), .C(n426), .Q(n421) );
  OAI212 U545 ( .A(n421), .B(n764), .C(n765), .Q(n56) );
  INV2 U546 ( .A(n171), .Q(n794) );
  NAND22 U547 ( .A(B[22]), .B(A[22]), .Q(n127) );
  NOR23 U548 ( .A(B[15]), .B(A[15]), .Q(n185) );
  OAI210 U549 ( .A(n177), .B(n173), .C(n174), .Q(n432) );
  NAND22 U551 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NOR24 U552 ( .A(n113), .B(n151), .Q(n111) );
  NAND22 U553 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND22 U554 ( .A(n766), .B(n71), .Q(n10) );
  NOR24 U555 ( .A(A[27]), .B(B[27]), .Q(n79) );
  NOR22 U557 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND22 U558 ( .A(n111), .B(n84), .Q(n82) );
  INV1 U559 ( .A(n268), .Q(n812) );
  INV0 U560 ( .A(n145), .Q(n787) );
  INV2 U561 ( .A(n73), .Q(n769) );
  NOR22 U562 ( .A(A[16]), .B(B[16]), .Q(n176) );
  INV1 U563 ( .A(n432), .Q(n795) );
  NAND21 U564 ( .A(n799), .B(n190), .Q(n188) );
  NAND21 U565 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND21 U566 ( .A(A[31]), .B(B[31]), .Q(n40) );
  XNR20 U567 ( .A(n34), .B(n812), .Q(SUM[4]) );
  CLKIN0 U568 ( .A(n239), .Q(n821) );
  INV0 U569 ( .A(n266), .Q(n815) );
  NOR20 U570 ( .A(n194), .B(n806), .Q(n190) );
  INV0 U571 ( .A(n231), .Q(n801) );
  INV0 U572 ( .A(n265), .Q(n814) );
  INV0 U573 ( .A(n255), .Q(n818) );
  NAND20 U574 ( .A(n811), .B(n272), .Q(n35) );
  NOR22 U575 ( .A(B[8]), .B(A[8]), .Q(n244) );
  INV2 U576 ( .A(n39), .Q(n759) );
  NAND20 U577 ( .A(n814), .B(n266), .Q(n34) );
  NAND20 U578 ( .A(n816), .B(n261), .Q(n33) );
  NAND22 U579 ( .A(n769), .B(n797), .Q(n596) );
  INV3 U580 ( .A(n219), .Q(n799) );
  INV3 U581 ( .A(n504), .Q(n819) );
  INV3 U582 ( .A(n82), .Q(n775) );
  NAND22 U583 ( .A(n258), .B(n250), .Q(n248) );
  NOR21 U584 ( .A(n271), .B(n274), .Q(n269) );
  NAND20 U585 ( .A(n239), .B(n800), .Q(n226) );
  AOI211 U586 ( .A(n504), .B(n800), .C(n801), .Q(n227) );
  NAND22 U587 ( .A(n799), .B(n810), .Q(n208) );
  AOI210 U588 ( .A(n796), .B(n810), .C(n809), .Q(n209) );
  INV3 U589 ( .A(n213), .Q(n809) );
  AOI210 U590 ( .A(n796), .B(n190), .C(n191), .Q(n189) );
  AOI211 U591 ( .A(n432), .B(n792), .C(n791), .Q(n159) );
  AOI210 U592 ( .A(n789), .B(n122), .C(n123), .Q(n121) );
  INV3 U593 ( .A(n420), .Q(n807) );
  NOR21 U594 ( .A(n260), .B(n265), .Q(n258) );
  INV3 U595 ( .A(n51), .Q(n761) );
  INV3 U596 ( .A(n230), .Q(n800) );
  INV3 U597 ( .A(n212), .Q(n810) );
  INV3 U598 ( .A(n185), .Q(n802) );
  INV3 U599 ( .A(n107), .Q(n777) );
  INV3 U600 ( .A(n70), .Q(n766) );
  INV0 U601 ( .A(n88), .Q(n781) );
  INV0 U602 ( .A(n126), .Q(n783) );
  INV0 U603 ( .A(n194), .Q(n804) );
  INV3 U604 ( .A(n244), .Q(n822) );
  NAND22 U605 ( .A(n817), .B(n253), .Q(n31) );
  INV3 U606 ( .A(n252), .Q(n817) );
  INV3 U607 ( .A(n117), .Q(n772) );
  INV3 U608 ( .A(n223), .Q(n798) );
  INV3 U609 ( .A(n173), .Q(n793) );
  INV3 U610 ( .A(n176), .Q(n808) );
  INV3 U611 ( .A(n195), .Q(n803) );
  INV3 U612 ( .A(n271), .Q(n811) );
  INV3 U613 ( .A(n260), .Q(n816) );
  INV3 U614 ( .A(n274), .Q(n823) );
  INV3 U615 ( .A(n277), .Q(n825) );
  INV3 U616 ( .A(n278), .Q(n827) );
  NOR21 U617 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NAND22 U618 ( .A(A[4]), .B(B[4]), .Q(n266) );
  INV3 U619 ( .A(n50), .Q(n760) );
  NOR21 U620 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U621 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U622 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U623 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NOR21 U624 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U625 ( .A(A[0]), .B(B[0]), .Q(n281) );
  INV3 U626 ( .A(n280), .Q(n826) );
  NOR21 U627 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U628 ( .A(n818), .B(n256), .Q(n32) );
  XNR21 U629 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XOR20 U630 ( .A(n758), .B(n22), .Q(SUM[16]) );
  NAND20 U631 ( .A(n808), .B(n177), .Q(n22) );
  NAND20 U632 ( .A(n100), .B(n782), .Q(n13) );
  NAND20 U633 ( .A(n762), .B(n62), .Q(n9) );
  NAND22 U634 ( .A(n759), .B(n40), .Q(n7) );
  XNR21 U635 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NAND20 U636 ( .A(n174), .B(n793), .Q(n21) );
  NAND20 U637 ( .A(n778), .B(n107), .Q(n14) );
  XNR21 U638 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND20 U639 ( .A(n788), .B(n145), .Q(n18) );
  XNR21 U640 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U641 ( .A(n156), .B(n756), .Q(n19) );
  XNR21 U642 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND20 U643 ( .A(n753), .B(n792), .Q(n20) );
  NAND20 U644 ( .A(n785), .B(n138), .Q(n17) );
  NAND20 U645 ( .A(n772), .B(n118), .Q(n15) );
  NAND20 U646 ( .A(n783), .B(n127), .Q(n16) );
  XNR21 U647 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U648 ( .A(n820), .B(n242), .Q(n29) );
  XNR21 U649 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U650 ( .A(n800), .B(n231), .Q(n28) );
  NAND20 U651 ( .A(n798), .B(n224), .Q(n27) );
  XNR21 U652 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U653 ( .A(n810), .B(n213), .Q(n26) );
  XNR21 U654 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U655 ( .A(n206), .B(n805), .Q(n25) );
  XNR21 U656 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U657 ( .A(n804), .B(n195), .Q(n24) );
  XNR21 U658 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U659 ( .A(n802), .B(n186), .Q(n23) );
  XOR20 U660 ( .A(n30), .B(n813), .Q(SUM[8]) );
  NAND20 U661 ( .A(n822), .B(n245), .Q(n30) );
  XOR21 U662 ( .A(n33), .B(n262), .Q(SUM[5]) );
  XOR21 U663 ( .A(n36), .B(n825), .Q(SUM[2]) );
  NAND22 U664 ( .A(n823), .B(n275), .Q(n36) );
  XNR21 U665 ( .A(n35), .B(n273), .Q(SUM[3]) );
  INV3 U666 ( .A(n38), .Q(SUM[0]) );
  NAND22 U667 ( .A(n826), .B(n281), .Q(n38) );
  XOR21 U668 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U669 ( .A(n827), .B(n279), .Q(n37) );
  NAND22 U670 ( .A(n111), .B(n44), .Q(n42) );
  NAND22 U671 ( .A(n111), .B(n97), .Q(n91) );
  CLKIN0 U672 ( .A(n137), .Q(n785) );
endmodule


module adder_22 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_22_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_21_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n50,
         n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n77, n78, n80, n81, n82, n83, n84, n85,
         n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103, n106,
         n107, n108, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n126, n127, n128, n129, n130, n135, n136,
         n137, n138, n139, n140, n141, n144, n145, n146, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n162, n163, n164, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n191, n194, n195, n196, n197,
         n198, n204, n205, n206, n207, n208, n209, n212, n213, n214, n219,
         n220, n221, n222, n224, n225, n226, n227, n230, n231, n232, n239,
         n240, n241, n242, n243, n244, n245, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n265, n266, n268, n269, n270, n271, n272, n273, n274, n275, n277,
         n278, n279, n280, n281, n420, n429, n430, n433, n434, n436, n437,
         n506, n507, n508, n581, n582, n584, n586, n587, n593, n594, n596,
         n600, n601, n602, n671, n678, n759, n760, n763, n764, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n920,
         n921, n922;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U65 ( .A(n82), .B(n845), .C(n83), .Q(n81) );
  OAI212 U77 ( .A(n91), .B(n845), .C(n92), .Q(n90) );
  OAI212 U141 ( .A(n140), .B(n845), .C(n141), .Q(n139) );
  OAI212 U165 ( .A(n158), .B(n845), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n885), .B(n845), .C(n882), .Q(n164) );
  OAI212 U197 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U219 ( .A(n197), .B(n904), .C(n198), .Q(n196) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U257 ( .A(n226), .B(n904), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n915), .B(n904), .C(n913), .Q(n232) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U329 ( .A(n274), .B(n921), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U495 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U476 ( .A(n73), .B(n845), .C(n74), .Q(n72) );
  OAI212 U505 ( .A(n862), .B(n845), .C(n857), .Q(n108) );
  OAI212 U395 ( .A(n129), .B(n845), .C(n130), .Q(n128) );
  OAI212 U404 ( .A(n120), .B(n845), .C(n121), .Q(n119) );
  OAI212 U426 ( .A(n151), .B(n845), .C(n671), .Q(n146) );
  OAI212 U436 ( .A(n89), .B(n436), .C(n80), .Q(n78) );
  OAI212 U440 ( .A(n244), .B(n904), .C(n245), .Q(n243) );
  OAI212 U441 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U449 ( .A(n53), .B(n845), .C(n54), .Q(n52) );
  OAI212 U502 ( .A(n760), .B(n878), .C(n89), .Q(n85) );
  AOI212 U356 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U451 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U465 ( .A(n113), .B(n671), .C(n114), .Q(n112) );
  OAI212 U488 ( .A(n176), .B(n845), .C(n177), .Q(n175) );
  OAI212 U408 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U422 ( .A(n42), .B(n845), .C(n43), .Q(n41) );
  OAI212 U469 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U491 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U517 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  CLKIN3 U349 ( .A(n155), .Q(n871) );
  NAND21 U350 ( .A(n860), .B(n118), .Q(n15) );
  NOR22 U351 ( .A(B[13]), .B(A[13]), .Q(n841) );
  NOR23 U352 ( .A(B[13]), .B(A[13]), .Q(n205) );
  OAI211 U353 ( .A(n194), .B(n901), .C(n195), .Q(n191) );
  AOI212 U354 ( .A(n183), .B(n204), .C(n184), .Q(n182) );
  NAND28 U355 ( .A(n600), .B(n114), .Q(n508) );
  NAND28 U357 ( .A(n861), .B(n872), .Q(n600) );
  NOR23 U358 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR24 U359 ( .A(B[12]), .B(A[12]), .Q(n212) );
  INV8 U360 ( .A(n212), .Q(n899) );
  OAI212 U361 ( .A(n126), .B(n866), .C(n127), .Q(n123) );
  NOR22 U362 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NAND20 U363 ( .A(n876), .B(n100), .Q(n13) );
  NOR23 U364 ( .A(n70), .B(n6), .Q(n66) );
  NOR22 U365 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR23 U366 ( .A(n194), .B(n586), .Q(n183) );
  NOR22 U367 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND22 U368 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND24 U369 ( .A(n429), .B(n430), .Q(SUM[27]) );
  NOR21 U370 ( .A(n436), .B(n88), .Q(n77) );
  NAND22 U371 ( .A(n97), .B(n77), .Q(n6) );
  NOR22 U372 ( .A(n155), .B(n162), .Q(n153) );
  INV3 U373 ( .A(n151), .Q(n874) );
  BUF6 U374 ( .A(n99), .Q(n844) );
  NOR21 U375 ( .A(n113), .B(n151), .Q(n111) );
  NAND22 U376 ( .A(n183), .B(n898), .Q(n181) );
  INV8 U377 ( .A(n596), .Q(n898) );
  NAND24 U378 ( .A(n907), .B(n899), .Q(n596) );
  NOR21 U379 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR21 U380 ( .A(n850), .B(n6), .Q(n55) );
  INV3 U381 ( .A(n507), .Q(n843) );
  INV3 U382 ( .A(n175), .Q(n889) );
  NAND22 U383 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NAND23 U384 ( .A(A[9]), .B(B[9]), .Q(n242) );
  AOI211 U385 ( .A(n890), .B(n897), .C(n191), .Q(n189) );
  NAND22 U386 ( .A(n897), .B(n888), .Q(n188) );
  XOR21 U387 ( .A(n33), .B(n262), .Q(SUM[5]) );
  XOR21 U388 ( .A(n32), .B(n257), .Q(SUM[6]) );
  XNR21 U389 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XNR21 U390 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XNR21 U391 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND23 U392 ( .A(n888), .B(n899), .Q(n208) );
  NAND22 U393 ( .A(n763), .B(n764), .Q(SUM[14]) );
  OAI212 U394 ( .A(n213), .B(n841), .C(n206), .Q(n204) );
  OAI210 U396 ( .A(n213), .B(n841), .C(n206), .Q(n420) );
  BUF2 U397 ( .A(n587), .Q(n842) );
  INV6 U398 ( .A(n152), .Q(n872) );
  NOR21 U399 ( .A(n126), .B(n865), .Q(n122) );
  NAND21 U400 ( .A(n871), .B(n156), .Q(n19) );
  NOR20 U401 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NOR22 U402 ( .A(n117), .B(n126), .Q(n115) );
  NOR22 U403 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR21 U405 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR21 U406 ( .A(B[8]), .B(A[8]), .Q(n244) );
  INV3 U407 ( .A(n135), .Q(n865) );
  NOR21 U409 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NAND21 U410 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NOR24 U411 ( .A(B[11]), .B(A[11]), .Q(n587) );
  NAND22 U412 ( .A(A[11]), .B(B[11]), .Q(n224) );
  OAI212 U413 ( .A(n188), .B(n904), .C(n189), .Q(n187) );
  NAND26 U414 ( .A(n135), .B(n115), .Q(n113) );
  AOI210 U415 ( .A(n872), .B(n135), .C(n136), .Q(n130) );
  AOI210 U416 ( .A(n872), .B(n122), .C(n123), .Q(n121) );
  NOR23 U417 ( .A(n587), .B(n230), .Q(n221) );
  INV1 U418 ( .A(n194), .Q(n906) );
  OAI212 U419 ( .A(n64), .B(n845), .C(n65), .Q(n63) );
  AOI212 U420 ( .A(n112), .B(n84), .C(n85), .Q(n83) );
  NAND21 U421 ( .A(A[21]), .B(B[21]), .Q(n138) );
  CLKIN0 U423 ( .A(n842), .Q(n909) );
  NAND21 U424 ( .A(n886), .B(n231), .Q(n28) );
  INV0 U425 ( .A(n231), .Q(n891) );
  OAI212 U427 ( .A(n127), .B(n437), .C(n118), .Q(n116) );
  NOR21 U428 ( .A(B[23]), .B(A[23]), .Q(n437) );
  OAI212 U429 ( .A(n102), .B(n845), .C(n103), .Q(n101) );
  CLKIN6 U430 ( .A(n153), .Q(n873) );
  NAND26 U431 ( .A(n506), .B(n174), .Q(n172) );
  NAND24 U432 ( .A(n895), .B(n884), .Q(n506) );
  CLKIN3 U433 ( .A(n437), .Q(n860) );
  NAND28 U434 ( .A(n889), .B(n883), .Q(n594) );
  XOR22 U435 ( .A(n22), .B(n845), .Q(SUM[16]) );
  INV1 U437 ( .A(n230), .Q(n886) );
  NAND20 U438 ( .A(n884), .B(n174), .Q(n21) );
  NAND28 U439 ( .A(n593), .B(n594), .Q(SUM[17]) );
  NAND21 U442 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND28 U443 ( .A(n581), .B(n582), .Q(SUM[19]) );
  NAND28 U444 ( .A(n879), .B(n870), .Q(n582) );
  NOR22 U445 ( .A(n181), .B(n219), .Q(n179) );
  INV6 U446 ( .A(n205), .Q(n907) );
  NOR22 U447 ( .A(A[25]), .B(B[25]), .Q(n99) );
  NOR21 U448 ( .A(B[7]), .B(A[7]), .Q(n252) );
  XNR22 U450 ( .A(n843), .B(n164), .Q(SUM[18]) );
  INV6 U452 ( .A(n172), .Q(n882) );
  XNR22 U453 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND22 U454 ( .A(n906), .B(n898), .Q(n584) );
  NAND22 U455 ( .A(n157), .B(n19), .Q(n581) );
  NAND24 U456 ( .A(n853), .B(n859), .Q(n430) );
  NOR22 U457 ( .A(n678), .B(n154), .Q(n671) );
  NOR24 U458 ( .A(n882), .B(n873), .Q(n678) );
  CLKIN2 U459 ( .A(n5), .Q(n856) );
  NAND21 U460 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NOR20 U461 ( .A(n271), .B(n274), .Q(n269) );
  OAI210 U462 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  NOR24 U463 ( .A(n678), .B(n154), .Q(n152) );
  AOI212 U464 ( .A(n508), .B(n893), .C(n894), .Q(n103) );
  NOR21 U466 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NOR21 U467 ( .A(B[5]), .B(A[5]), .Q(n260) );
  XNR22 U468 ( .A(n9), .B(n63), .Q(SUM[29]) );
  OAI212 U470 ( .A(n208), .B(n904), .C(n209), .Q(n207) );
  AOI210 U471 ( .A(n890), .B(n899), .C(n900), .Q(n209) );
  INV3 U472 ( .A(n220), .Q(n890) );
  XNR22 U473 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NOR21 U474 ( .A(B[26]), .B(A[26]), .Q(n760) );
  INV1 U475 ( .A(n97), .Q(n877) );
  OAI211 U477 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  AOI210 U478 ( .A(n508), .B(n44), .C(n45), .Q(n43) );
  NAND21 U479 ( .A(n863), .B(n127), .Q(n16) );
  OAI212 U480 ( .A(n107), .B(n844), .C(n100), .Q(n98) );
  NAND21 U481 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND22 U482 ( .A(A[10]), .B(B[10]), .Q(n231) );
  XNR22 U483 ( .A(n15), .B(n119), .Q(SUM[23]) );
  OAI212 U484 ( .A(n231), .B(n587), .C(n224), .Q(n222) );
  NOR22 U485 ( .A(B[10]), .B(A[10]), .Q(n230) );
  AOI211 U486 ( .A(n890), .B(n898), .C(n420), .Q(n198) );
  NAND20 U487 ( .A(n899), .B(n213), .Q(n26) );
  NOR21 U489 ( .A(B[15]), .B(A[15]), .Q(n185) );
  XNR22 U490 ( .A(n10), .B(n72), .Q(SUM[28]) );
  INV2 U492 ( .A(n113), .Q(n861) );
  AOI211 U493 ( .A(n240), .B(n886), .C(n891), .Q(n227) );
  NAND21 U494 ( .A(A[17]), .B(B[17]), .Q(n174) );
  XNR22 U496 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND22 U497 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND22 U498 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U499 ( .A(n893), .B(n107), .Q(n14) );
  INV1 U500 ( .A(n107), .Q(n894) );
  AOI211 U501 ( .A(n508), .B(n855), .C(n856), .Q(n74) );
  CLKIN6 U503 ( .A(n157), .Q(n879) );
  NAND23 U504 ( .A(n171), .B(n153), .Q(n151) );
  NAND22 U506 ( .A(n874), .B(n135), .Q(n129) );
  NAND22 U507 ( .A(n874), .B(n122), .Q(n120) );
  XNR22 U508 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U509 ( .A(n25), .B(n207), .Q(SUM[13]) );
  CLKIN3 U510 ( .A(n136), .Q(n866) );
  XNR22 U511 ( .A(n8), .B(n52), .Q(SUM[30]) );
  INV0 U512 ( .A(n126), .Q(n863) );
  AOI212 U513 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NAND24 U514 ( .A(A[12]), .B(B[12]), .Q(n213) );
  INV3 U515 ( .A(n173), .Q(n884) );
  NOR22 U516 ( .A(B[16]), .B(A[16]), .Q(n176) );
  XNR22 U518 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NOR24 U519 ( .A(n113), .B(n151), .Q(n602) );
  CLKIN3 U520 ( .A(n508), .Q(n857) );
  AOI211 U521 ( .A(n508), .B(n97), .C(n98), .Q(n92) );
  XNR22 U522 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NOR22 U523 ( .A(B[21]), .B(A[21]), .Q(n601) );
  AOI211 U524 ( .A(n872), .B(n867), .C(n868), .Q(n141) );
  NAND21 U525 ( .A(n602), .B(n893), .Q(n102) );
  NAND22 U526 ( .A(n602), .B(n855), .Q(n73) );
  NAND21 U527 ( .A(n602), .B(n55), .Q(n53) );
  CLKIN2 U528 ( .A(n602), .Q(n862) );
  OAI212 U529 ( .A(n185), .B(n195), .C(n186), .Q(n184) );
  NAND22 U530 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NOR22 U531 ( .A(B[15]), .B(A[15]), .Q(n586) );
  AOI211 U532 ( .A(n508), .B(n66), .C(n67), .Q(n65) );
  NAND21 U533 ( .A(n906), .B(n195), .Q(n24) );
  NOR22 U534 ( .A(B[19]), .B(A[19]), .Q(n155) );
  INV2 U535 ( .A(n601), .Q(n864) );
  NOR22 U536 ( .A(n601), .B(n144), .Q(n135) );
  NAND24 U537 ( .A(n433), .B(n434), .Q(SUM[25]) );
  NOR23 U538 ( .A(B[27]), .B(A[27]), .Q(n436) );
  NAND21 U539 ( .A(n111), .B(n97), .Q(n91) );
  NAND20 U540 ( .A(n914), .B(n242), .Q(n29) );
  BUF15 U541 ( .A(n178), .Q(n845) );
  INV0 U542 ( .A(n61), .Q(n849) );
  INV1 U543 ( .A(n106), .Q(n893) );
  CLKIN3 U544 ( .A(n196), .Q(n887) );
  NAND20 U545 ( .A(n867), .B(n145), .Q(n18) );
  NAND20 U546 ( .A(n896), .B(n177), .Q(n22) );
  NAND22 U547 ( .A(n849), .B(n62), .Q(n9) );
  NAND22 U548 ( .A(n852), .B(n71), .Q(n10) );
  INV0 U549 ( .A(n70), .Q(n852) );
  NAND22 U550 ( .A(n918), .B(n245), .Q(n30) );
  INV2 U551 ( .A(n244), .Q(n918) );
  INV1 U552 ( .A(n51), .Q(n847) );
  NAND22 U553 ( .A(n24), .B(n196), .Q(n763) );
  INV0 U554 ( .A(n171), .Q(n885) );
  NAND20 U555 ( .A(n907), .B(n206), .Q(n25) );
  NAND20 U556 ( .A(n171), .B(n881), .Q(n158) );
  AOI210 U557 ( .A(n172), .B(n881), .C(n880), .Q(n159) );
  NAND20 U558 ( .A(n888), .B(n898), .Q(n197) );
  NOR20 U559 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND20 U560 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND21 U561 ( .A(n602), .B(n66), .Q(n64) );
  NOR20 U562 ( .A(B[18]), .B(A[18]), .Q(n759) );
  NOR20 U563 ( .A(n46), .B(n6), .Q(n44) );
  CLKIN3 U564 ( .A(n60), .Q(n851) );
  AOI210 U565 ( .A(n112), .B(n55), .C(n56), .Q(n54) );
  NAND20 U566 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U567 ( .A(n239), .B(n886), .Q(n226) );
  INV2 U568 ( .A(n241), .Q(n914) );
  AOI210 U569 ( .A(n60), .B(n848), .C(n847), .Q(n47) );
  NOR22 U570 ( .A(n844), .B(n106), .Q(n97) );
  NAND20 U571 ( .A(n59), .B(n848), .Q(n46) );
  INV2 U572 ( .A(n265), .Q(n911) );
  NOR20 U573 ( .A(n241), .B(n244), .Q(n239) );
  NOR20 U574 ( .A(n260), .B(n265), .Q(n258) );
  NOR20 U575 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR20 U576 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR20 U577 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND20 U578 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U579 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U580 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND20 U581 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U582 ( .A(n175), .B(n21), .Q(n593) );
  INV3 U583 ( .A(n21), .Q(n883) );
  NAND22 U584 ( .A(n905), .B(n887), .Q(n764) );
  INV3 U585 ( .A(n24), .Q(n905) );
  INV3 U586 ( .A(n19), .Q(n870) );
  NAND22 U587 ( .A(n874), .B(n867), .Q(n140) );
  INV3 U588 ( .A(n584), .Q(n897) );
  NAND22 U589 ( .A(n892), .B(n186), .Q(n23) );
  INV3 U590 ( .A(n586), .Q(n892) );
  INV3 U591 ( .A(n176), .Q(n896) );
  NAND22 U592 ( .A(n864), .B(n138), .Q(n17) );
  NOR21 U593 ( .A(n173), .B(n176), .Q(n171) );
  NOR21 U594 ( .A(n759), .B(n880), .Q(n507) );
  INV3 U595 ( .A(n759), .Q(n881) );
  XNR21 U596 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND22 U597 ( .A(n909), .B(n224), .Q(n27) );
  INV3 U598 ( .A(n213), .Q(n900) );
  INV3 U599 ( .A(n204), .Q(n901) );
  INV3 U600 ( .A(n145), .Q(n868) );
  INV3 U601 ( .A(n177), .Q(n895) );
  NAND20 U602 ( .A(n602), .B(n44), .Q(n42) );
  INV3 U603 ( .A(n144), .Q(n867) );
  INV3 U604 ( .A(n163), .Q(n880) );
  INV3 U605 ( .A(n219), .Q(n888) );
  INV3 U606 ( .A(n239), .Q(n915) );
  NAND22 U607 ( .A(n875), .B(n858), .Q(n434) );
  NAND21 U608 ( .A(n13), .B(n101), .Q(n433) );
  INV3 U609 ( .A(n13), .Q(n875) );
  NAND21 U610 ( .A(n11), .B(n81), .Q(n429) );
  INV3 U611 ( .A(n11), .Q(n853) );
  INV3 U612 ( .A(n101), .Q(n858) );
  INV3 U613 ( .A(n81), .Q(n859) );
  INV3 U614 ( .A(n6), .Q(n855) );
  INV0 U615 ( .A(n240), .Q(n913) );
  INV3 U616 ( .A(n59), .Q(n850) );
  AOI211 U617 ( .A(n903), .B(n258), .C(n259), .Q(n257) );
  NAND20 U618 ( .A(n239), .B(n221), .Q(n219) );
  INV3 U619 ( .A(n247), .Q(n904) );
  INV3 U620 ( .A(n268), .Q(n903) );
  INV3 U621 ( .A(n277), .Q(n921) );
  AOI211 U622 ( .A(n903), .B(n911), .C(n910), .Q(n262) );
  NAND22 U623 ( .A(n912), .B(n261), .Q(n33) );
  INV3 U624 ( .A(n266), .Q(n910) );
  XOR21 U625 ( .A(n30), .B(n904), .Q(SUM[8]) );
  NAND22 U626 ( .A(n908), .B(n256), .Q(n32) );
  INV3 U627 ( .A(n255), .Q(n908) );
  NAND22 U628 ( .A(n869), .B(n89), .Q(n12) );
  INV3 U629 ( .A(n760), .Q(n869) );
  NAND22 U630 ( .A(n848), .B(n51), .Q(n8) );
  XNR21 U631 ( .A(n34), .B(n903), .Q(SUM[4]) );
  NAND22 U632 ( .A(n911), .B(n266), .Q(n34) );
  NAND22 U633 ( .A(n917), .B(n253), .Q(n31) );
  INV3 U634 ( .A(n252), .Q(n917) );
  XNR21 U635 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U636 ( .A(n902), .B(n272), .Q(n35) );
  INV3 U637 ( .A(n271), .Q(n902) );
  NOR21 U638 ( .A(n61), .B(n70), .Q(n59) );
  INV3 U639 ( .A(n844), .Q(n876) );
  NAND22 U640 ( .A(n854), .B(n80), .Q(n11) );
  INV3 U641 ( .A(n436), .Q(n854) );
  NAND22 U642 ( .A(n111), .B(n84), .Q(n82) );
  NOR22 U643 ( .A(n760), .B(n877), .Q(n84) );
  XNR21 U644 ( .A(n29), .B(n243), .Q(SUM[9]) );
  INV1 U645 ( .A(n98), .Q(n878) );
  INV3 U646 ( .A(n260), .Q(n912) );
  XOR21 U647 ( .A(n36), .B(n921), .Q(SUM[2]) );
  NAND22 U648 ( .A(n916), .B(n275), .Q(n36) );
  INV3 U649 ( .A(n274), .Q(n916) );
  AOI211 U650 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NAND22 U651 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U652 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U653 ( .A(n252), .B(n255), .Q(n250) );
  XOR21 U654 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U655 ( .A(n922), .B(n279), .Q(n37) );
  INV3 U656 ( .A(n278), .Q(n922) );
  XNR21 U657 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U658 ( .A(n846), .B(n40), .Q(n7) );
  NAND20 U659 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR20 U660 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV3 U661 ( .A(n50), .Q(n848) );
  NOR20 U662 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND20 U663 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U664 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NOR20 U665 ( .A(B[2]), .B(A[2]), .Q(n274) );
  INV3 U666 ( .A(n39), .Q(n846) );
  NAND20 U667 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND20 U668 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND20 U669 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U670 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND20 U671 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND20 U672 ( .A(A[7]), .B(B[7]), .Q(n253) );
  INV3 U673 ( .A(n38), .Q(SUM[0]) );
  NAND22 U674 ( .A(n920), .B(n281), .Q(n38) );
  INV3 U675 ( .A(n280), .Q(n920) );
  NOR20 U676 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U677 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NOR20 U678 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND20 U679 ( .A(A[1]), .B(B[1]), .Q(n279) );
  OAI210 U680 ( .A(n219), .B(n904), .C(n220), .Q(n214) );
  OAI210 U681 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI210 U682 ( .A(n850), .B(n5), .C(n851), .Q(n56) );
  NOR21 U683 ( .A(B[24]), .B(A[24]), .Q(n106) );
endmodule


module adder_21 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_21_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_20_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n418, n486, n560,
         n567, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780;

  OAI212 U51 ( .A(n73), .B(n718), .C(n74), .Q(n72) );
  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U65 ( .A(n82), .B(n718), .C(n83), .Q(n81) );
  OAI212 U105 ( .A(n152), .B(n113), .C(n114), .Q(n112) );
  OAI212 U135 ( .A(n145), .B(n717), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n718), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n718), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n757), .B(n718), .C(n758), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  AOI212 U249 ( .A(n221), .B(n240), .C(n222), .Q(n220) );
  OAI212 U275 ( .A(n241), .B(n245), .C(n242), .Q(n240) );
  AOI212 U290 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n721), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U403 ( .A(n255), .B(n715), .C(n710), .Q(n254) );
  OAI212 U389 ( .A(n113), .B(n152), .C(n114), .Q(n418) );
  OAI212 U349 ( .A(n197), .B(n722), .C(n198), .Q(n196) );
  OAI212 U427 ( .A(n774), .B(n722), .C(n772), .Q(n232) );
  OAI212 U452 ( .A(n188), .B(n722), .C(n189), .Q(n187) );
  OAI212 U477 ( .A(n226), .B(n722), .C(n227), .Q(n225) );
  XNR22 U484 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI212 U510 ( .A(n208), .B(n722), .C(n209), .Q(n207) );
  OAI212 U371 ( .A(n248), .B(n268), .C(n249), .Q(n560) );
  OAI212 U390 ( .A(n266), .B(n260), .C(n261), .Q(n486) );
  OAI212 U465 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  XNR22 U414 ( .A(n13), .B(n101), .Q(SUM[25]) );
  OAI212 U493 ( .A(n176), .B(n718), .C(n177), .Q(n175) );
  OAI212 U350 ( .A(n42), .B(n718), .C(n43), .Q(n41) );
  OAI212 U392 ( .A(n126), .B(n748), .C(n127), .Q(n123) );
  OAI212 U415 ( .A(n102), .B(n718), .C(n103), .Q(n101) );
  OAI212 U446 ( .A(n744), .B(n718), .C(n743), .Q(n108) );
  OAI212 U474 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U481 ( .A(n88), .B(n739), .C(n89), .Q(n85) );
  OAI212 U485 ( .A(n730), .B(n5), .C(n731), .Q(n56) );
  OAI212 U516 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U521 ( .A(n64), .B(n718), .C(n65), .Q(n63) );
  NAND22 U351 ( .A(A[19]), .B(B[19]), .Q(n156) );
  INV3 U352 ( .A(n152), .Q(n753) );
  NOR24 U353 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR23 U354 ( .A(n244), .B(n713), .Q(n239) );
  INV1 U355 ( .A(n212), .Q(n766) );
  XNR22 U356 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NOR22 U357 ( .A(B[23]), .B(A[23]), .Q(n117) );
  XNR22 U358 ( .A(n26), .B(n214), .Q(SUM[12]) );
  XNR22 U359 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND23 U360 ( .A(n97), .B(n77), .Q(n6) );
  NOR21 U361 ( .A(n730), .B(n6), .Q(n55) );
  INV3 U362 ( .A(n712), .Q(n713) );
  NOR21 U363 ( .A(n61), .B(n70), .Q(n59) );
  AOI211 U364 ( .A(n418), .B(n84), .C(n85), .Q(n83) );
  NOR21 U365 ( .A(n70), .B(n6), .Q(n66) );
  NOR23 U366 ( .A(n205), .B(n212), .Q(n203) );
  AOI211 U367 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  INV3 U368 ( .A(n213), .Q(n765) );
  INV3 U369 ( .A(n256), .Q(n709) );
  OAI212 U370 ( .A(n194), .B(n764), .C(n195), .Q(n191) );
  NAND21 U372 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NAND22 U373 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND22 U374 ( .A(n752), .B(n122), .Q(n120) );
  INV3 U375 ( .A(n135), .Q(n747) );
  INV3 U376 ( .A(n709), .Q(n710) );
  NAND22 U377 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND23 U378 ( .A(n203), .B(n183), .Q(n181) );
  OAI212 U379 ( .A(n244), .B(n722), .C(n245), .Q(n243) );
  INV6 U380 ( .A(n560), .Q(n722) );
  INV3 U381 ( .A(n767), .Q(n711) );
  INV3 U382 ( .A(n241), .Q(n712) );
  NOR21 U383 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR22 U384 ( .A(A[12]), .B(B[12]), .Q(n212) );
  NAND21 U385 ( .A(n769), .B(n203), .Q(n197) );
  INV2 U386 ( .A(n219), .Q(n769) );
  OAI212 U387 ( .A(n120), .B(n718), .C(n121), .Q(n119) );
  INV2 U388 ( .A(n203), .Q(n763) );
  NAND20 U391 ( .A(n776), .B(n253), .Q(n31) );
  CLKIN0 U393 ( .A(n244), .Q(n775) );
  CLKIN0 U394 ( .A(n713), .Q(n773) );
  NOR23 U395 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND22 U396 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NOR23 U397 ( .A(n181), .B(n219), .Q(n179) );
  AOI210 U398 ( .A(n418), .B(n55), .C(n56), .Q(n54) );
  AOI210 U399 ( .A(n418), .B(n734), .C(n735), .Q(n74) );
  NOR22 U400 ( .A(B[26]), .B(A[26]), .Q(n88) );
  INV2 U401 ( .A(n220), .Q(n767) );
  NOR23 U402 ( .A(n252), .B(n255), .Q(n250) );
  AOI212 U404 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  OAI212 U405 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  INV0 U406 ( .A(n239), .Q(n774) );
  OAI211 U407 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NAND21 U408 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND21 U409 ( .A(n751), .B(n156), .Q(n19) );
  AOI211 U410 ( .A(n112), .B(n97), .C(n98), .Q(n92) );
  OAI211 U411 ( .A(n53), .B(n718), .C(n54), .Q(n52) );
  NOR22 U412 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND20 U413 ( .A(A[21]), .B(B[21]), .Q(n138) );
  INV1 U416 ( .A(n204), .Q(n764) );
  AOI211 U417 ( .A(n767), .B(n203), .C(n204), .Q(n198) );
  NAND21 U418 ( .A(n769), .B(n766), .Q(n208) );
  XNR22 U419 ( .A(n9), .B(n63), .Q(SUM[29]) );
  INV0 U420 ( .A(n205), .Q(n762) );
  AOI212 U421 ( .A(n767), .B(n190), .C(n191), .Q(n189) );
  NAND22 U422 ( .A(A[16]), .B(B[16]), .Q(n177) );
  OAI211 U423 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  NAND20 U424 ( .A(n761), .B(n195), .Q(n24) );
  NOR22 U425 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND21 U426 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR21 U428 ( .A(n173), .B(n176), .Q(n171) );
  OAI211 U429 ( .A(n129), .B(n718), .C(n130), .Q(n128) );
  NOR22 U430 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR24 U431 ( .A(A[7]), .B(B[7]), .Q(n252) );
  NAND21 U432 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NOR24 U433 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NOR23 U434 ( .A(A[14]), .B(B[14]), .Q(n194) );
  XOR21 U435 ( .A(n30), .B(n722), .Q(SUM[8]) );
  XNR22 U436 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XOR22 U437 ( .A(n22), .B(n718), .Q(SUM[16]) );
  CLKBU15 U438 ( .A(n178), .Q(n718) );
  OAI212 U439 ( .A(n151), .B(n718), .C(n152), .Q(n146) );
  OAI212 U440 ( .A(n91), .B(n718), .C(n92), .Q(n90) );
  NOR21 U441 ( .A(n194), .B(n763), .Q(n190) );
  XNR22 U442 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND23 U443 ( .A(n135), .B(n115), .Q(n113) );
  NOR22 U444 ( .A(n117), .B(n126), .Q(n115) );
  NOR22 U445 ( .A(n717), .B(n144), .Q(n135) );
  NOR24 U447 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NAND21 U448 ( .A(n261), .B(n778), .Q(n33) );
  XOR22 U449 ( .A(n33), .B(n262), .Q(SUM[5]) );
  XNR22 U450 ( .A(n29), .B(n243), .Q(SUM[9]) );
  XNR22 U451 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XOR21 U453 ( .A(n32), .B(n715), .Q(SUM[6]) );
  AOI212 U454 ( .A(n716), .B(n258), .C(n486), .Q(n715) );
  NOR21 U455 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR23 U456 ( .A(B[9]), .B(A[9]), .Q(n241) );
  XNR22 U457 ( .A(n24), .B(n196), .Q(SUM[14]) );
  XNR22 U458 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NOR21 U459 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NAND20 U460 ( .A(n111), .B(n55), .Q(n53) );
  XNR22 U461 ( .A(n18), .B(n146), .Q(SUM[20]) );
  AOI211 U462 ( .A(n714), .B(n770), .C(n771), .Q(n227) );
  INV1 U463 ( .A(n230), .Q(n770) );
  XNR22 U464 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND21 U466 ( .A(n111), .B(n97), .Q(n91) );
  NOR21 U467 ( .A(B[27]), .B(A[27]), .Q(n79) );
  OAI211 U468 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NAND21 U469 ( .A(A[26]), .B(B[26]), .Q(n89) );
  XNR22 U470 ( .A(n139), .B(n17), .Q(SUM[21]) );
  XNR22 U471 ( .A(n15), .B(n119), .Q(SUM[23]) );
  XNR22 U472 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND21 U473 ( .A(B[13]), .B(A[13]), .Q(n206) );
  XNR22 U475 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NAND23 U476 ( .A(n567), .B(n253), .Q(n251) );
  NAND21 U478 ( .A(A[7]), .B(B[7]), .Q(n253) );
  OAI210 U479 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI211 U480 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  AOI211 U482 ( .A(n753), .B(n122), .C(n123), .Q(n121) );
  NOR24 U483 ( .A(n185), .B(n194), .Q(n183) );
  INV2 U486 ( .A(n772), .Q(n714) );
  NAND21 U487 ( .A(A[9]), .B(B[9]), .Q(n242) );
  INV1 U488 ( .A(n240), .Q(n772) );
  NOR23 U489 ( .A(n223), .B(n230), .Q(n221) );
  NAND20 U490 ( .A(n239), .B(n770), .Q(n226) );
  XNR22 U491 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND21 U492 ( .A(A[15]), .B(B[15]), .Q(n186) );
  OAI211 U494 ( .A(n219), .B(n722), .C(n711), .Q(n214) );
  NAND24 U495 ( .A(n239), .B(n221), .Q(n219) );
  CLKIN6 U496 ( .A(n252), .Q(n776) );
  OAI212 U497 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  NAND21 U498 ( .A(n770), .B(n231), .Q(n28) );
  NAND22 U499 ( .A(A[10]), .B(B[10]), .Q(n231) );
  XNR22 U500 ( .A(n20), .B(n164), .Q(SUM[18]) );
  OAI212 U501 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  NAND21 U502 ( .A(n766), .B(n213), .Q(n26) );
  NAND22 U503 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NOR22 U504 ( .A(n79), .B(n88), .Q(n77) );
  INV0 U505 ( .A(n79), .Q(n733) );
  INV3 U506 ( .A(n151), .Q(n752) );
  NOR23 U507 ( .A(n113), .B(n151), .Q(n111) );
  NAND20 U508 ( .A(n752), .B(n135), .Q(n129) );
  INV1 U509 ( .A(n144), .Q(n750) );
  NAND21 U511 ( .A(A[24]), .B(B[24]), .Q(n107) );
  AOI210 U512 ( .A(n753), .B(n135), .C(n136), .Q(n130) );
  NOR21 U513 ( .A(n99), .B(n106), .Q(n97) );
  CLKIN0 U514 ( .A(n106), .Q(n741) );
  NOR22 U515 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NAND21 U517 ( .A(n111), .B(n741), .Q(n102) );
  NAND21 U518 ( .A(n190), .B(n769), .Q(n188) );
  INV1 U519 ( .A(n5), .Q(n735) );
  NAND20 U520 ( .A(n737), .B(n100), .Q(n13) );
  NAND22 U522 ( .A(n732), .B(n71), .Q(n10) );
  INV0 U523 ( .A(n70), .Q(n732) );
  INV0 U524 ( .A(n162), .Q(n754) );
  INV2 U525 ( .A(n271), .Q(n725) );
  NOR20 U526 ( .A(n271), .B(n274), .Q(n269) );
  INV1 U527 ( .A(n6), .Q(n734) );
  NAND21 U528 ( .A(n111), .B(n66), .Q(n64) );
  INV3 U529 ( .A(n268), .Q(n716) );
  CLKIN3 U530 ( .A(n60), .Q(n731) );
  CLKIN3 U531 ( .A(n59), .Q(n730) );
  NAND20 U532 ( .A(n171), .B(n754), .Q(n158) );
  CLKIN0 U533 ( .A(n171), .Q(n757) );
  NAND20 U534 ( .A(n775), .B(n245), .Q(n30) );
  INV0 U535 ( .A(n99), .Q(n737) );
  AOI210 U536 ( .A(n418), .B(n66), .C(n67), .Q(n65) );
  INV0 U537 ( .A(n136), .Q(n748) );
  INV0 U538 ( .A(n61), .Q(n729) );
  INV0 U539 ( .A(n717), .Q(n746) );
  NAND22 U540 ( .A(n138), .B(n746), .Q(n17) );
  NAND20 U541 ( .A(n745), .B(n127), .Q(n16) );
  NAND20 U542 ( .A(n742), .B(n118), .Q(n15) );
  AOI210 U543 ( .A(n60), .B(n728), .C(n727), .Q(n47) );
  NAND20 U544 ( .A(n777), .B(n710), .Q(n32) );
  INV0 U545 ( .A(n255), .Q(n777) );
  NAND20 U546 ( .A(n779), .B(n266), .Q(n34) );
  NAND20 U547 ( .A(n59), .B(n728), .Q(n46) );
  INV0 U548 ( .A(n223), .Q(n768) );
  INV2 U549 ( .A(n265), .Q(n779) );
  INV0 U550 ( .A(n266), .Q(n780) );
  NOR20 U551 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NAND20 U552 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U553 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND20 U554 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND22 U555 ( .A(n111), .B(n734), .Q(n73) );
  INV3 U556 ( .A(n111), .Q(n744) );
  NAND20 U557 ( .A(n111), .B(n44), .Q(n42) );
  NAND22 U558 ( .A(n171), .B(n153), .Q(n151) );
  NOR20 U559 ( .A(n46), .B(n6), .Q(n44) );
  NAND22 U560 ( .A(n111), .B(n84), .Q(n82) );
  NAND22 U561 ( .A(n752), .B(n750), .Q(n140) );
  NAND22 U562 ( .A(n258), .B(n250), .Q(n248) );
  INV3 U563 ( .A(n277), .Q(n721) );
  NAND22 U564 ( .A(n759), .B(n177), .Q(n22) );
  CLKIN0 U565 ( .A(n176), .Q(n759) );
  XNR21 U566 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND22 U567 ( .A(n736), .B(n89), .Q(n12) );
  INV3 U568 ( .A(n88), .Q(n736) );
  XNR21 U569 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND22 U570 ( .A(n741), .B(n107), .Q(n14) );
  INV3 U571 ( .A(n112), .Q(n743) );
  INV3 U572 ( .A(n126), .Q(n745) );
  INV0 U573 ( .A(n117), .Q(n742) );
  NAND22 U574 ( .A(n728), .B(n51), .Q(n8) );
  XNR21 U575 ( .A(n34), .B(n716), .Q(SUM[4]) );
  XNR21 U576 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U577 ( .A(n725), .B(n272), .Q(n35) );
  NAND22 U578 ( .A(n733), .B(n80), .Q(n11) );
  NAND22 U579 ( .A(n729), .B(n62), .Q(n9) );
  INV3 U580 ( .A(n231), .Q(n771) );
  NAND20 U581 ( .A(n750), .B(n145), .Q(n18) );
  NAND22 U582 ( .A(n760), .B(n186), .Q(n23) );
  INV3 U583 ( .A(n185), .Q(n760) );
  NAND20 U584 ( .A(n773), .B(n242), .Q(n29) );
  NAND20 U585 ( .A(n768), .B(n224), .Q(n27) );
  NAND20 U586 ( .A(n762), .B(n206), .Q(n25) );
  NAND22 U587 ( .A(n754), .B(n163), .Q(n20) );
  INV0 U588 ( .A(n172), .Q(n758) );
  INV0 U589 ( .A(n155), .Q(n751) );
  NOR21 U590 ( .A(n126), .B(n747), .Q(n122) );
  AOI211 U591 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NOR22 U592 ( .A(n155), .B(n162), .Q(n153) );
  NAND22 U593 ( .A(n709), .B(n776), .Q(n567) );
  AOI211 U594 ( .A(n716), .B(n779), .C(n780), .Q(n262) );
  INV0 U595 ( .A(n260), .Q(n778) );
  NOR21 U596 ( .A(n88), .B(n738), .Q(n84) );
  INV2 U597 ( .A(n97), .Q(n738) );
  AOI210 U598 ( .A(n172), .B(n754), .C(n755), .Q(n159) );
  INV3 U599 ( .A(n163), .Q(n755) );
  AOI211 U600 ( .A(n112), .B(n741), .C(n740), .Q(n103) );
  INV3 U601 ( .A(n107), .Q(n740) );
  AOI211 U602 ( .A(n753), .B(n750), .C(n749), .Q(n141) );
  INV0 U603 ( .A(n145), .Q(n749) );
  INV0 U604 ( .A(n98), .Q(n739) );
  AOI210 U605 ( .A(n418), .B(n44), .C(n45), .Q(n43) );
  INV3 U606 ( .A(n51), .Q(n727) );
  AOI211 U607 ( .A(n767), .B(n766), .C(n765), .Q(n209) );
  INV0 U608 ( .A(n173), .Q(n756) );
  NAND20 U609 ( .A(n756), .B(n174), .Q(n21) );
  XOR21 U610 ( .A(n36), .B(n721), .Q(SUM[2]) );
  NAND22 U611 ( .A(n724), .B(n275), .Q(n36) );
  INV3 U612 ( .A(n274), .Q(n724) );
  XOR21 U613 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U614 ( .A(n723), .B(n279), .Q(n37) );
  INV3 U615 ( .A(n278), .Q(n723) );
  NOR21 U616 ( .A(B[18]), .B(A[18]), .Q(n162) );
  XNR21 U617 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U618 ( .A(n726), .B(n40), .Q(n7) );
  NAND20 U619 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND22 U620 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND22 U621 ( .A(B[8]), .B(A[8]), .Q(n245) );
  NAND20 U622 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND22 U623 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND20 U624 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND20 U625 ( .A(A[28]), .B(B[28]), .Q(n71) );
  BUF6 U626 ( .A(n137), .Q(n717) );
  INV3 U627 ( .A(n50), .Q(n728) );
  NOR20 U628 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U629 ( .A(n39), .Q(n726) );
  NOR20 U630 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND20 U631 ( .A(A[3]), .B(B[3]), .Q(n272) );
  INV3 U632 ( .A(n38), .Q(SUM[0]) );
  NAND22 U633 ( .A(n720), .B(n281), .Q(n38) );
  INV3 U634 ( .A(n280), .Q(n720) );
  NOR20 U635 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NOR20 U636 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND20 U637 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U638 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NOR20 U639 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND20 U640 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NOR23 U641 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR22 U642 ( .A(A[17]), .B(B[17]), .Q(n173) );
  NOR20 U643 ( .A(n260), .B(n265), .Q(n258) );
  NOR22 U644 ( .A(B[19]), .B(A[19]), .Q(n155) );
  INV1 U645 ( .A(n194), .Q(n761) );
  NOR21 U646 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR22 U647 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR22 U648 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U649 ( .A(B[20]), .B(A[20]), .Q(n144) );
endmodule


module adder_20 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_20_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_19_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n191, n194, n195, n196,
         n197, n198, n203, n204, n205, n206, n207, n208, n209, n212, n213,
         n214, n219, n220, n221, n222, n223, n224, n225, n226, n227, n230,
         n231, n232, n239, n240, n241, n242, n243, n244, n245, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n265, n266, n268, n269, n270, n271, n272, n273,
         n274, n275, n277, n278, n279, n280, n281, n421, n423, n426, n430,
         n498, n500, n501, n503, n509, n510, n577, n581, n582, n585, n589,
         n590, n593, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n814;

  OAI212 U165 ( .A(n158), .B(n743), .C(n159), .Q(n157) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U227 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U563 ( .A(n274), .B(n811), .C(n275), .Q(n273) );
  OAI212 U500 ( .A(n510), .B(n46), .C(n47), .Q(n45) );
  OAI212 U518 ( .A(n42), .B(n740), .C(n43), .Q(n41) );
  OAI212 U519 ( .A(n99), .B(n107), .C(n100), .Q(n98) );
  OAI212 U409 ( .A(n793), .B(n743), .C(n791), .Q(n164) );
  OAI212 U466 ( .A(n761), .B(n743), .C(n759), .Q(n108) );
  AOI212 U509 ( .A(n172), .B(n153), .C(n498), .Q(n500) );
  OAI212 U511 ( .A(n82), .B(n740), .C(n83), .Q(n81) );
  OAI212 U538 ( .A(n223), .B(n231), .C(n224), .Q(n222) );
  OAI212 U442 ( .A(n241), .B(n245), .C(n242), .Q(n240) );
  OAI212 U479 ( .A(n64), .B(n740), .C(n65), .Q(n63) );
  OAI212 U514 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U529 ( .A(n53), .B(n740), .C(n54), .Q(n52) );
  OAI212 U530 ( .A(n107), .B(n99), .C(n100), .Q(n430) );
  AOI212 U546 ( .A(n77), .B(n430), .C(n78), .Q(n510) );
  OAI212 U551 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U481 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U573 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  INV0 U349 ( .A(n780), .Q(n738) );
  INV3 U350 ( .A(n220), .Q(n780) );
  NAND22 U351 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND21 U352 ( .A(A[7]), .B(B[7]), .Q(n253) );
  INV2 U353 ( .A(n194), .Q(n789) );
  INV2 U354 ( .A(n742), .Q(n759) );
  NOR24 U355 ( .A(A[25]), .B(B[25]), .Q(n99) );
  NOR22 U356 ( .A(n88), .B(n764), .Q(n84) );
  NOR24 U357 ( .A(n162), .B(n155), .Q(n153) );
  INV2 U358 ( .A(n173), .Q(n792) );
  NAND20 U359 ( .A(n171), .B(n779), .Q(n158) );
  NOR23 U360 ( .A(n230), .B(n223), .Q(n221) );
  INV2 U361 ( .A(n163), .Q(n777) );
  NAND24 U362 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NOR24 U363 ( .A(B[18]), .B(A[18]), .Q(n162) );
  INV15 U364 ( .A(n781), .Q(n740) );
  AOI212 U365 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR23 U366 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR24 U367 ( .A(n194), .B(n185), .Q(n183) );
  NOR24 U368 ( .A(B[15]), .B(A[15]), .Q(n185) );
  AOI211 U369 ( .A(n503), .B(n97), .C(n430), .Q(n92) );
  OAI211 U370 ( .A(n500), .B(n113), .C(n114), .Q(n503) );
  NAND28 U371 ( .A(n97), .B(n77), .Q(n6) );
  NOR23 U372 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NAND26 U373 ( .A(n593), .B(n74), .Q(n72) );
  NOR23 U374 ( .A(n99), .B(n106), .Q(n97) );
  OAI212 U375 ( .A(n743), .B(n91), .C(n92), .Q(n90) );
  NAND21 U376 ( .A(B[27]), .B(A[27]), .Q(n80) );
  NOR23 U377 ( .A(n205), .B(n212), .Q(n203) );
  NOR22 U378 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR24 U379 ( .A(n79), .B(n88), .Q(n77) );
  NAND26 U380 ( .A(n509), .B(n80), .Q(n78) );
  INV0 U381 ( .A(n88), .Q(n758) );
  NAND21 U382 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NOR24 U383 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR23 U384 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR23 U385 ( .A(n61), .B(n70), .Q(n59) );
  NOR23 U386 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND23 U387 ( .A(n59), .B(n746), .Q(n46) );
  CLKIN3 U388 ( .A(n135), .Q(n770) );
  NAND24 U389 ( .A(n153), .B(n171), .Q(n151) );
  NOR22 U390 ( .A(n271), .B(n274), .Q(n269) );
  NOR21 U391 ( .A(n260), .B(n265), .Q(n258) );
  NAND24 U392 ( .A(n203), .B(n183), .Q(n181) );
  NAND22 U393 ( .A(A[24]), .B(B[24]), .Q(n107) );
  INV3 U394 ( .A(n268), .Q(n804) );
  NAND22 U395 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND23 U396 ( .A(B[16]), .B(A[16]), .Q(n177) );
  NOR23 U397 ( .A(n252), .B(n255), .Q(n250) );
  AOI212 U398 ( .A(n772), .B(n501), .C(n771), .Q(n577) );
  INV3 U399 ( .A(n774), .Q(n739) );
  CLKIN3 U400 ( .A(n247), .Q(n802) );
  OAI212 U401 ( .A(n129), .B(n743), .C(n130), .Q(n128) );
  NAND22 U402 ( .A(A[25]), .B(B[25]), .Q(n100) );
  INV3 U403 ( .A(n510), .Q(n753) );
  CLKIN15 U404 ( .A(n741), .Q(n742) );
  NAND22 U405 ( .A(n44), .B(n111), .Q(n42) );
  NOR22 U406 ( .A(n46), .B(n6), .Q(n44) );
  NAND21 U407 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NAND22 U408 ( .A(A[3]), .B(B[3]), .Q(n272) );
  CLKIN0 U410 ( .A(n205), .Q(n790) );
  NOR23 U411 ( .A(n70), .B(n6), .Q(n66) );
  CLKIN2 U412 ( .A(n231), .Q(n797) );
  INV3 U413 ( .A(n97), .Q(n764) );
  NOR23 U414 ( .A(n173), .B(n176), .Q(n171) );
  AOI210 U415 ( .A(n780), .B(n203), .C(n204), .Q(n198) );
  CLKIN6 U416 ( .A(n79), .Q(n754) );
  NOR24 U417 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR23 U418 ( .A(n241), .B(n244), .Q(n239) );
  INV0 U419 ( .A(n241), .Q(n801) );
  NOR23 U420 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND21 U421 ( .A(n746), .B(n51), .Q(n8) );
  NOR22 U422 ( .A(n117), .B(n126), .Q(n423) );
  INV0 U423 ( .A(n117), .Q(n760) );
  NAND28 U424 ( .A(n135), .B(n115), .Q(n113) );
  CLKIN15 U425 ( .A(n743), .Q(n781) );
  CLKIN0 U426 ( .A(n223), .Q(n783) );
  AOI212 U427 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  INV0 U428 ( .A(n252), .Q(n803) );
  AOI211 U429 ( .A(n774), .B(n769), .C(n767), .Q(n141) );
  INV6 U430 ( .A(n112), .Q(n741) );
  OAI210 U431 ( .A(n245), .B(n241), .C(n242), .Q(n421) );
  NOR24 U432 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NAND22 U433 ( .A(n776), .B(n769), .Q(n140) );
  OAI212 U434 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  NOR24 U435 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND21 U436 ( .A(n111), .B(n84), .Q(n82) );
  CLKIN3 U437 ( .A(n171), .Q(n793) );
  INV2 U438 ( .A(n111), .Q(n761) );
  NAND22 U439 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND22 U440 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NOR22 U441 ( .A(B[24]), .B(A[24]), .Q(n106) );
  CLKBU15 U443 ( .A(n178), .Q(n743) );
  NAND21 U444 ( .A(A[13]), .B(B[13]), .Q(n206) );
  AOI211 U445 ( .A(n135), .B(n774), .C(n501), .Q(n130) );
  NAND21 U446 ( .A(n789), .B(n203), .Q(n426) );
  XNR22 U447 ( .A(n7), .B(n41), .Q(SUM[31]) );
  INV0 U448 ( .A(n137), .Q(n773) );
  OAI211 U449 ( .A(n145), .B(n137), .C(n138), .Q(n501) );
  AOI212 U450 ( .A(n742), .B(n84), .C(n85), .Q(n83) );
  NAND21 U451 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NOR24 U452 ( .A(B[29]), .B(A[29]), .Q(n61) );
  INV6 U453 ( .A(n50), .Q(n746) );
  NOR24 U454 ( .A(B[30]), .B(A[30]), .Q(n50) );
  AOI211 U455 ( .A(n774), .B(n122), .C(n768), .Q(n121) );
  INV4 U456 ( .A(n500), .Q(n774) );
  INV4 U457 ( .A(n6), .Q(n756) );
  AOI212 U458 ( .A(n742), .B(n55), .C(n56), .Q(n54) );
  NAND22 U459 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NOR23 U460 ( .A(n117), .B(n126), .Q(n115) );
  NOR24 U461 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR22 U462 ( .A(B[10]), .B(A[10]), .Q(n230) );
  INV2 U463 ( .A(n219), .Q(n784) );
  NOR24 U464 ( .A(n181), .B(n219), .Q(n179) );
  NAND22 U465 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND24 U467 ( .A(n239), .B(n221), .Q(n219) );
  NOR24 U468 ( .A(B[9]), .B(A[9]), .Q(n241) );
  CLKIN1 U469 ( .A(n162), .Q(n779) );
  INV1 U470 ( .A(n106), .Q(n765) );
  OAI211 U471 ( .A(n151), .B(n743), .C(n739), .Q(n146) );
  XNR22 U472 ( .A(n9), .B(n63), .Q(SUM[29]) );
  OAI212 U473 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  AOI212 U474 ( .A(n60), .B(n746), .C(n745), .Q(n47) );
  NAND21 U475 ( .A(A[1]), .B(B[1]), .Q(n279) );
  XOR21 U476 ( .A(n30), .B(n802), .Q(SUM[8]) );
  NOR24 U477 ( .A(n144), .B(n137), .Q(n135) );
  NAND21 U478 ( .A(n776), .B(n122), .Q(n120) );
  NAND22 U480 ( .A(A[12]), .B(B[12]), .Q(n213) );
  OAI211 U482 ( .A(n88), .B(n762), .C(n89), .Q(n85) );
  INV3 U483 ( .A(n98), .Q(n762) );
  AOI212 U484 ( .A(n742), .B(n765), .C(n766), .Q(n103) );
  NAND24 U485 ( .A(n589), .B(n590), .Q(SUM[28]) );
  NAND24 U486 ( .A(n750), .B(n752), .Q(n590) );
  CLKIN6 U487 ( .A(n72), .Q(n752) );
  OAI212 U488 ( .A(n5), .B(n748), .C(n749), .Q(n56) );
  OAI212 U489 ( .A(n5), .B(n70), .C(n71), .Q(n67) );
  NAND21 U490 ( .A(n111), .B(n97), .Q(n91) );
  NOR24 U491 ( .A(B[17]), .B(A[17]), .Q(n173) );
  AOI212 U492 ( .A(n742), .B(n66), .C(n67), .Q(n65) );
  XNR22 U493 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XNR22 U494 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NAND24 U495 ( .A(n755), .B(n781), .Q(n593) );
  NAND20 U496 ( .A(n769), .B(n145), .Q(n18) );
  INV0 U497 ( .A(n145), .Q(n767) );
  NAND23 U498 ( .A(A[20]), .B(B[20]), .Q(n145) );
  AOI210 U499 ( .A(n585), .B(n779), .C(n777), .Q(n159) );
  NAND22 U501 ( .A(n55), .B(n111), .Q(n53) );
  NOR22 U502 ( .A(n748), .B(n6), .Q(n55) );
  NAND21 U503 ( .A(n765), .B(n107), .Q(n14) );
  AOI212 U504 ( .A(n742), .B(n756), .C(n753), .Q(n74) );
  NOR24 U505 ( .A(B[19]), .B(A[19]), .Q(n155) );
  OAI211 U506 ( .A(n120), .B(n743), .C(n121), .Q(n119) );
  OAI211 U507 ( .A(n140), .B(n743), .C(n141), .Q(n139) );
  NAND22 U508 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND22 U510 ( .A(A[14]), .B(B[14]), .Q(n195) );
  OAI212 U512 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  NAND21 U513 ( .A(n111), .B(n765), .Q(n102) );
  NAND22 U515 ( .A(n111), .B(n66), .Q(n64) );
  NOR24 U516 ( .A(n151), .B(n113), .Q(n111) );
  NAND21 U517 ( .A(n787), .B(n213), .Q(n26) );
  INV1 U520 ( .A(n213), .Q(n785) );
  AOI212 U521 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  INV2 U522 ( .A(n204), .Q(n786) );
  NOR24 U523 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND20 U524 ( .A(n784), .B(n203), .Q(n197) );
  NAND20 U525 ( .A(n789), .B(n195), .Q(n24) );
  AOI212 U526 ( .A(n742), .B(n44), .C(n45), .Q(n43) );
  OAI211 U527 ( .A(n188), .B(n802), .C(n189), .Q(n187) );
  OAI211 U528 ( .A(n197), .B(n802), .C(n198), .Q(n196) );
  OAI211 U531 ( .A(n208), .B(n802), .C(n209), .Q(n207) );
  OAI211 U532 ( .A(n226), .B(n802), .C(n227), .Q(n225) );
  OAI211 U533 ( .A(n799), .B(n802), .C(n800), .Q(n232) );
  OAI212 U534 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND20 U535 ( .A(n747), .B(n62), .Q(n9) );
  NOR24 U536 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND22 U537 ( .A(A[26]), .B(B[26]), .Q(n89) );
  OAI211 U539 ( .A(n219), .B(n802), .C(n738), .Q(n214) );
  XNR22 U540 ( .A(n13), .B(n101), .Q(SUM[25]) );
  OAI212 U541 ( .A(n102), .B(n740), .C(n103), .Q(n101) );
  AOI212 U542 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  NAND21 U543 ( .A(n776), .B(n135), .Q(n129) );
  INV0 U544 ( .A(n185), .Q(n795) );
  NOR24 U545 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR23 U547 ( .A(B[20]), .B(A[20]), .Q(n144) );
  OAI212 U548 ( .A(n155), .B(n163), .C(n156), .Q(n154) );
  OAI212 U549 ( .A(n155), .B(n163), .C(n156), .Q(n498) );
  INV2 U550 ( .A(n155), .Q(n775) );
  AOI212 U552 ( .A(n136), .B(n423), .C(n116), .Q(n114) );
  OAI211 U553 ( .A(n244), .B(n802), .C(n245), .Q(n243) );
  NOR22 U554 ( .A(B[8]), .B(A[8]), .Q(n244) );
  INV3 U555 ( .A(n59), .Q(n748) );
  AOI212 U556 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  AOI212 U557 ( .A(n153), .B(n585), .C(n154), .Q(n152) );
  AOI210 U558 ( .A(n780), .B(n787), .C(n785), .Q(n209) );
  NAND21 U559 ( .A(B[23]), .B(A[23]), .Q(n118) );
  OAI212 U560 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U561 ( .A(n177), .B(n173), .C(n174), .Q(n585) );
  NAND22 U562 ( .A(A[22]), .B(B[22]), .Q(n127) );
  OAI211 U564 ( .A(n176), .B(n743), .C(n177), .Q(n175) );
  OAI211 U565 ( .A(n194), .B(n786), .C(n195), .Q(n191) );
  NAND22 U566 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND22 U567 ( .A(n794), .B(n177), .Q(n22) );
  NAND21 U568 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV1 U569 ( .A(n20), .Q(n778) );
  CLKIN0 U570 ( .A(n239), .Q(n799) );
  CLKIN2 U571 ( .A(n172), .Q(n791) );
  AOI211 U572 ( .A(n804), .B(n258), .C(n259), .Q(n257) );
  CLKIN1 U574 ( .A(n421), .Q(n800) );
  INV0 U575 ( .A(n212), .Q(n787) );
  INV0 U576 ( .A(n230), .Q(n796) );
  NAND21 U577 ( .A(n20), .B(n164), .Q(n581) );
  CLKIN3 U578 ( .A(n10), .Q(n750) );
  CLKIN3 U579 ( .A(n164), .Q(n782) );
  INV0 U580 ( .A(n266), .Q(n809) );
  NAND20 U581 ( .A(n779), .B(n163), .Q(n20) );
  INV0 U582 ( .A(n265), .Q(n808) );
  INV0 U583 ( .A(n244), .Q(n798) );
  INV0 U584 ( .A(n278), .Q(n812) );
  INV0 U585 ( .A(n274), .Q(n810) );
  INV0 U586 ( .A(n271), .Q(n805) );
  NOR22 U587 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND21 U588 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND21 U589 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U590 ( .A(n39), .Q(n744) );
  NAND21 U591 ( .A(n100), .B(n763), .Q(n13) );
  NAND20 U592 ( .A(n810), .B(n275), .Q(n36) );
  NAND20 U593 ( .A(n805), .B(n272), .Q(n35) );
  INV3 U594 ( .A(n151), .Q(n776) );
  INV3 U595 ( .A(n73), .Q(n755) );
  NAND22 U596 ( .A(n111), .B(n756), .Q(n73) );
  NAND20 U597 ( .A(n784), .B(n788), .Q(n188) );
  AOI211 U598 ( .A(n780), .B(n788), .C(n191), .Q(n189) );
  INV3 U599 ( .A(n426), .Q(n788) );
  NAND22 U600 ( .A(n778), .B(n782), .Q(n582) );
  NAND22 U601 ( .A(n258), .B(n250), .Q(n248) );
  NOR21 U602 ( .A(n126), .B(n770), .Q(n122) );
  NAND20 U603 ( .A(n239), .B(n796), .Q(n226) );
  AOI211 U604 ( .A(n421), .B(n796), .C(n797), .Q(n227) );
  NAND20 U605 ( .A(n784), .B(n787), .Q(n208) );
  AOI210 U606 ( .A(n804), .B(n808), .C(n809), .Q(n262) );
  INV3 U607 ( .A(n51), .Q(n745) );
  NAND22 U608 ( .A(n751), .B(n71), .Q(n10) );
  INV3 U609 ( .A(n70), .Q(n751) );
  NAND22 U610 ( .A(n757), .B(n754), .Q(n509) );
  INV3 U611 ( .A(n89), .Q(n757) );
  INV3 U612 ( .A(n144), .Q(n769) );
  INV0 U613 ( .A(n277), .Q(n811) );
  INV3 U614 ( .A(n126), .Q(n772) );
  INV3 U615 ( .A(n260), .Q(n807) );
  INV3 U616 ( .A(n255), .Q(n806) );
  INV3 U617 ( .A(n61), .Q(n747) );
  INV3 U618 ( .A(n176), .Q(n794) );
  CLKIN3 U619 ( .A(n577), .Q(n768) );
  INV3 U620 ( .A(n127), .Q(n771) );
  NOR21 U621 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U622 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV3 U623 ( .A(n107), .Q(n766) );
  NOR21 U624 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U625 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U626 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND22 U627 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NOR21 U628 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U629 ( .A(n280), .Q(n814) );
  NOR21 U630 ( .A(B[0]), .B(A[0]), .Q(n280) );
  XOR21 U631 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND20 U632 ( .A(n807), .B(n261), .Q(n33) );
  NAND22 U633 ( .A(n744), .B(n40), .Q(n7) );
  NAND21 U634 ( .A(n10), .B(n72), .Q(n589) );
  XOR20 U635 ( .A(n743), .B(n22), .Q(SUM[16]) );
  XNR21 U636 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U637 ( .A(n783), .B(n224), .Q(n27) );
  XNR21 U638 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U639 ( .A(n796), .B(n231), .Q(n28) );
  XNR21 U640 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U641 ( .A(n206), .B(n790), .Q(n25) );
  XNR21 U642 ( .A(n24), .B(n196), .Q(SUM[14]) );
  XNR21 U643 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U644 ( .A(n803), .B(n253), .Q(n31) );
  NAND20 U645 ( .A(n798), .B(n245), .Q(n30) );
  XOR21 U646 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND20 U647 ( .A(n812), .B(n279), .Q(n37) );
  XNR20 U648 ( .A(n34), .B(n804), .Q(SUM[4]) );
  NAND20 U649 ( .A(n808), .B(n266), .Q(n34) );
  NAND22 U650 ( .A(n581), .B(n582), .Q(SUM[18]) );
  XNR21 U651 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U652 ( .A(n242), .B(n801), .Q(n29) );
  XNR21 U653 ( .A(n26), .B(n214), .Q(SUM[12]) );
  XNR21 U654 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U655 ( .A(n795), .B(n186), .Q(n23) );
  XOR20 U656 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND20 U657 ( .A(n806), .B(n256), .Q(n32) );
  XNR21 U658 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XOR21 U659 ( .A(n36), .B(n811), .Q(SUM[2]) );
  XNR21 U660 ( .A(n12), .B(n90), .Q(SUM[26]) );
  XNR21 U661 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NAND20 U662 ( .A(n174), .B(n792), .Q(n21) );
  XNR21 U663 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND20 U664 ( .A(n127), .B(n772), .Q(n16) );
  XNR21 U665 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND20 U666 ( .A(n760), .B(n118), .Q(n15) );
  XNR21 U667 ( .A(n18), .B(n146), .Q(SUM[20]) );
  XNR21 U668 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR21 U669 ( .A(n17), .B(n139), .Q(SUM[21]) );
  NAND20 U670 ( .A(n773), .B(n138), .Q(n17) );
  XNR21 U671 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U672 ( .A(n156), .B(n775), .Q(n19) );
  INV3 U673 ( .A(n38), .Q(SUM[0]) );
  NAND22 U674 ( .A(n814), .B(n281), .Q(n38) );
  NAND20 U675 ( .A(n754), .B(n80), .Q(n11) );
  NAND22 U676 ( .A(n758), .B(n89), .Q(n12) );
  CLKIN0 U677 ( .A(n99), .Q(n763) );
  INV3 U678 ( .A(n60), .Q(n749) );
endmodule


module adder_19 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_19_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_18_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n55, n56, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n194, n195, n196,
         n197, n198, n204, n205, n206, n207, n208, n209, n212, n213, n214,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n230, n231,
         n232, n239, n240, n241, n242, n243, n244, n245, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n265, n266, n268, n269, n270, n272, n273, n274, n275,
         n277, n278, n279, n280, n281, n431, n432, n500, n503, n504, n507,
         n508, n511, n519, n521, n591, n592, n595, n596, n674, n675, n677,
         n682, n683, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U127 ( .A(n129), .B(n772), .C(n130), .Q(n128) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n772), .C(n141), .Q(n139) );
  OAI212 U159 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U165 ( .A(n158), .B(n772), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n803), .B(n772), .C(n799), .Q(n164) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n252), .B(n256), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n260), .B(n266), .C(n261), .Q(n259) );
  AOI212 U321 ( .A(n269), .B(n277), .C(n270), .Q(n268) );
  OAI212 U349 ( .A(n177), .B(n763), .C(n174), .Q(n172) );
  AOI212 U357 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  AOI212 U407 ( .A(n250), .B(n259), .C(n251), .Q(n249) );
  OAI212 U458 ( .A(n91), .B(n772), .C(n92), .Q(n90) );
  OAI212 U394 ( .A(n785), .B(n783), .C(n773), .Q(n232) );
  OAI212 U479 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U517 ( .A(n102), .B(n772), .C(n103), .Q(n101) );
  OAI212 U492 ( .A(n185), .B(n195), .C(n186), .Q(n184) );
  OAI212 U469 ( .A(n197), .B(n785), .C(n198), .Q(n196) );
  OAI212 U474 ( .A(n208), .B(n785), .C(n209), .Q(n207) );
  OAI212 U497 ( .A(n176), .B(n772), .C(n177), .Q(n511) );
  OAI212 U436 ( .A(n244), .B(n785), .C(n245), .Q(n243) );
  OAI212 U477 ( .A(n275), .B(n519), .C(n272), .Q(n270) );
  OAI212 U496 ( .A(n785), .B(n226), .C(n227), .Q(n225) );
  OAI212 U510 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U515 ( .A(n64), .B(n772), .C(n65), .Q(n63) );
  OAI212 U549 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U677 ( .A(n151), .B(n772), .C(n152), .Q(n146) );
  OAI212 U468 ( .A(n126), .B(n811), .C(n127), .Q(n123) );
  OAI212 U507 ( .A(n828), .B(n5), .C(n829), .Q(n56) );
  OAI212 U508 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U518 ( .A(n42), .B(n772), .C(n43), .Q(n41) );
  OAI212 U540 ( .A(n73), .B(n772), .C(n74), .Q(n72) );
  OAI212 U541 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND22 U350 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR23 U351 ( .A(A[13]), .B(B[13]), .Q(n205) );
  NOR22 U352 ( .A(n79), .B(n88), .Q(n77) );
  INV2 U353 ( .A(n252), .Q(n786) );
  INV8 U354 ( .A(n247), .Q(n785) );
  NOR21 U355 ( .A(n46), .B(n6), .Q(n44) );
  NAND23 U356 ( .A(n97), .B(n77), .Q(n6) );
  NOR23 U358 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR24 U359 ( .A(A[6]), .B(B[6]), .Q(n255) );
  NOR22 U360 ( .A(B[22]), .B(A[22]), .Q(n126) );
  AOI212 U361 ( .A(n761), .B(n84), .C(n85), .Q(n83) );
  NOR22 U362 ( .A(A[17]), .B(B[17]), .Q(n173) );
  CLKIN6 U363 ( .A(n762), .Q(n763) );
  AOI211 U364 ( .A(n761), .B(n832), .C(n831), .Q(n74) );
  CLKIN10 U365 ( .A(n759), .Q(n761) );
  AOI212 U366 ( .A(n800), .B(n122), .C(n123), .Q(n121) );
  INV2 U367 ( .A(n152), .Q(n800) );
  AOI211 U368 ( .A(n800), .B(n135), .C(n136), .Q(n130) );
  NOR23 U369 ( .A(A[9]), .B(B[9]), .Q(n241) );
  XNR22 U370 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U371 ( .A(n23), .B(n187), .Q(SUM[15]) );
  XNR22 U372 ( .A(n13), .B(n101), .Q(SUM[25]) );
  INV6 U373 ( .A(n112), .Q(n759) );
  INV4 U374 ( .A(n759), .Q(n760) );
  CLKIN4 U375 ( .A(n173), .Q(n762) );
  XOR22 U376 ( .A(n22), .B(n772), .Q(SUM[16]) );
  XOR22 U377 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NOR21 U378 ( .A(B[24]), .B(A[24]), .Q(n106) );
  CLKIN3 U379 ( .A(n511), .Q(n781) );
  NAND22 U380 ( .A(n806), .B(n777), .Q(n682) );
  XNR21 U381 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NOR22 U382 ( .A(n117), .B(n126), .Q(n115) );
  NOR23 U383 ( .A(n185), .B(n194), .Q(n183) );
  NOR22 U384 ( .A(n99), .B(n106), .Q(n97) );
  NOR21 U385 ( .A(B[28]), .B(A[28]), .Q(n70) );
  AOI211 U386 ( .A(n761), .B(n97), .C(n98), .Q(n92) );
  NOR21 U387 ( .A(n126), .B(n813), .Q(n122) );
  NOR22 U388 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND20 U389 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NOR23 U390 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND23 U391 ( .A(A[2]), .B(B[2]), .Q(n275) );
  INV3 U392 ( .A(n205), .Q(n826) );
  NAND24 U393 ( .A(n431), .B(n432), .Q(SUM[17]) );
  NAND23 U395 ( .A(n781), .B(n820), .Q(n432) );
  NAND24 U396 ( .A(n595), .B(n596), .Q(SUM[9]) );
  AOI211 U397 ( .A(n787), .B(n798), .C(n797), .Q(n262) );
  NAND28 U398 ( .A(n677), .B(n224), .Q(n222) );
  NAND20 U399 ( .A(A[21]), .B(B[21]), .Q(n138) );
  AOI211 U400 ( .A(n775), .B(n190), .C(n191), .Q(n189) );
  OAI211 U401 ( .A(n248), .B(n268), .C(n249), .Q(n764) );
  NAND22 U402 ( .A(B[3]), .B(A[3]), .Q(n272) );
  NAND20 U403 ( .A(n272), .B(n788), .Q(n35) );
  CLKIN0 U404 ( .A(n260), .Q(n793) );
  NOR23 U405 ( .A(n241), .B(n244), .Q(n239) );
  AOI212 U406 ( .A(n760), .B(n837), .C(n838), .Q(n103) );
  NOR24 U408 ( .A(n181), .B(n219), .Q(n179) );
  OAI212 U409 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  NOR21 U410 ( .A(B[1]), .B(A[1]), .Q(n278) );
  OAI211 U411 ( .A(n274), .B(n791), .C(n275), .Q(n273) );
  NOR22 U412 ( .A(n274), .B(n519), .Q(n269) );
  NAND23 U413 ( .A(B[8]), .B(A[8]), .Q(n245) );
  INV3 U414 ( .A(n519), .Q(n788) );
  OAI212 U415 ( .A(n805), .B(n772), .C(n801), .Q(n108) );
  NOR22 U416 ( .A(n260), .B(n265), .Q(n258) );
  NAND24 U417 ( .A(n809), .B(n779), .Q(n592) );
  CLKIN6 U418 ( .A(n119), .Q(n779) );
  NAND22 U419 ( .A(n848), .B(n780), .Q(n508) );
  NOR22 U420 ( .A(n255), .B(n252), .Q(n250) );
  XNR21 U421 ( .A(n34), .B(n787), .Q(SUM[4]) );
  NOR23 U422 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND22 U423 ( .A(n225), .B(n27), .Q(n767) );
  NAND28 U424 ( .A(n765), .B(n766), .Q(n768) );
  NAND28 U425 ( .A(n767), .B(n768), .Q(SUM[11]) );
  CLKIN6 U426 ( .A(n225), .Q(n765) );
  INV12 U427 ( .A(n27), .Q(n766) );
  NAND24 U428 ( .A(n507), .B(n508), .Q(SUM[22]) );
  NAND23 U429 ( .A(n250), .B(n258), .Q(n248) );
  NOR22 U430 ( .A(n763), .B(n176), .Q(n171) );
  NAND23 U431 ( .A(n171), .B(n153), .Q(n151) );
  AOI210 U432 ( .A(n761), .B(n66), .C(n67), .Q(n65) );
  AOI210 U433 ( .A(n683), .B(n823), .C(n822), .Q(n227) );
  CLKIN6 U434 ( .A(n157), .Q(n778) );
  NAND23 U435 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND24 U437 ( .A(n674), .B(n675), .Q(SUM[12]) );
  NAND22 U438 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND22 U439 ( .A(n157), .B(n19), .Q(n503) );
  OAI210 U440 ( .A(n245), .B(n241), .C(n242), .Q(n683) );
  NAND24 U441 ( .A(n795), .B(n774), .Q(n596) );
  NAND22 U442 ( .A(n243), .B(n29), .Q(n595) );
  CLKIN6 U443 ( .A(n243), .Q(n774) );
  OAI212 U444 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U445 ( .A(n188), .B(n785), .C(n189), .Q(n187) );
  NOR20 U446 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U447 ( .A(A[6]), .B(B[6]), .Q(n256) );
  INV6 U448 ( .A(n521), .Q(n825) );
  NAND24 U449 ( .A(n778), .B(n818), .Q(n504) );
  NAND20 U450 ( .A(n843), .B(n213), .Q(n26) );
  INV2 U451 ( .A(n136), .Q(n811) );
  INV3 U452 ( .A(n268), .Q(n787) );
  INV1 U453 ( .A(n265), .Q(n798) );
  NOR24 U454 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV1 U455 ( .A(n204), .Q(n824) );
  OAI212 U456 ( .A(n82), .B(n772), .C(n83), .Q(n81) );
  INV0 U457 ( .A(n244), .Q(n782) );
  NAND24 U459 ( .A(n822), .B(n816), .Q(n677) );
  CLKIN6 U460 ( .A(n223), .Q(n816) );
  XNR22 U461 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NOR23 U462 ( .A(n223), .B(n230), .Q(n221) );
  NAND24 U463 ( .A(n135), .B(n115), .Q(n113) );
  NAND22 U464 ( .A(A[4]), .B(B[4]), .Q(n266) );
  XNR22 U465 ( .A(n9), .B(n63), .Q(SUM[29]) );
  OAI212 U466 ( .A(n219), .B(n785), .C(n220), .Q(n214) );
  NAND22 U467 ( .A(A[24]), .B(B[24]), .Q(n107) );
  XNR22 U470 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND22 U471 ( .A(n111), .B(n837), .Q(n102) );
  NOR24 U472 ( .A(n113), .B(n151), .Q(n111) );
  INV1 U473 ( .A(n106), .Q(n837) );
  NOR24 U475 ( .A(n155), .B(n162), .Q(n153) );
  INV0 U476 ( .A(n155), .Q(n819) );
  NOR23 U478 ( .A(A[19]), .B(B[19]), .Q(n155) );
  NAND24 U480 ( .A(n826), .B(n843), .Q(n521) );
  NOR24 U481 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR24 U482 ( .A(B[11]), .B(A[11]), .Q(n223) );
  XNR22 U483 ( .A(n24), .B(n196), .Q(SUM[14]) );
  INV3 U484 ( .A(n220), .Q(n775) );
  NOR23 U485 ( .A(B[7]), .B(A[7]), .Q(n252) );
  CLKIN0 U486 ( .A(n763), .Q(n821) );
  OAI211 U487 ( .A(n176), .B(n772), .C(n177), .Q(n500) );
  NAND22 U488 ( .A(A[18]), .B(B[18]), .Q(n163) );
  INV3 U489 ( .A(n97), .Q(n836) );
  NAND22 U490 ( .A(n111), .B(n97), .Q(n91) );
  NOR23 U491 ( .A(n137), .B(n144), .Q(n135) );
  NAND24 U493 ( .A(n503), .B(n504), .Q(SUM[19]) );
  NOR22 U494 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NAND21 U495 ( .A(n16), .B(n128), .Q(n507) );
  CLKIN4 U498 ( .A(n128), .Q(n780) );
  NOR24 U499 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND21 U500 ( .A(B[17]), .B(A[17]), .Q(n174) );
  XNR22 U501 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND21 U502 ( .A(n804), .B(n122), .Q(n120) );
  NAND21 U503 ( .A(n214), .B(n26), .Q(n674) );
  XNR22 U504 ( .A(n31), .B(n254), .Q(SUM[7]) );
  INV6 U505 ( .A(n219), .Q(n784) );
  NAND26 U506 ( .A(n239), .B(n221), .Q(n219) );
  NAND21 U509 ( .A(A[26]), .B(B[26]), .Q(n89) );
  XNR22 U511 ( .A(n12), .B(n90), .Q(SUM[26]) );
  NAND21 U512 ( .A(A[15]), .B(B[15]), .Q(n186) );
  OAI210 U513 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  CLKIN1 U514 ( .A(n277), .Q(n791) );
  XNR22 U516 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND20 U519 ( .A(n239), .B(n823), .Q(n226) );
  INV1 U520 ( .A(n230), .Q(n823) );
  XNR22 U521 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND22 U522 ( .A(n784), .B(n190), .Q(n188) );
  NOR21 U523 ( .A(n194), .B(n521), .Q(n190) );
  INV1 U524 ( .A(n5), .Q(n831) );
  AOI212 U525 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI212 U526 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NAND21 U527 ( .A(n784), .B(n825), .Q(n197) );
  OAI211 U528 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NOR22 U529 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND21 U530 ( .A(B[19]), .B(A[19]), .Q(n156) );
  NAND26 U531 ( .A(n825), .B(n183), .Q(n181) );
  AOI212 U532 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  INV1 U533 ( .A(n772), .Q(n777) );
  NOR22 U534 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NAND22 U535 ( .A(B[12]), .B(A[12]), .Q(n213) );
  XNR22 U536 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NAND24 U537 ( .A(n591), .B(n592), .Q(SUM[23]) );
  XNR22 U538 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NOR24 U539 ( .A(A[3]), .B(B[3]), .Q(n519) );
  XNR22 U542 ( .A(n139), .B(n17), .Q(SUM[21]) );
  OAI212 U543 ( .A(n120), .B(n772), .C(n121), .Q(n119) );
  BUF15 U544 ( .A(n178), .Q(n772) );
  CLKIN3 U545 ( .A(n801), .Q(n770) );
  INV2 U546 ( .A(n761), .Q(n801) );
  NOR24 U547 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND22 U548 ( .A(n804), .B(n135), .Q(n129) );
  INV3 U550 ( .A(n151), .Q(n804) );
  NAND21 U551 ( .A(n111), .B(n84), .Q(n82) );
  NAND22 U552 ( .A(n111), .B(n66), .Q(n64) );
  NAND21 U553 ( .A(n111), .B(n44), .Q(n42) );
  NAND21 U554 ( .A(n111), .B(n55), .Q(n53) );
  NAND22 U555 ( .A(n111), .B(n832), .Q(n73) );
  INV2 U556 ( .A(n111), .Q(n805) );
  XOR22 U557 ( .A(n257), .B(n32), .Q(SUM[6]) );
  AOI212 U558 ( .A(n787), .B(n258), .C(n259), .Q(n257) );
  CLKIN0 U559 ( .A(n88), .Q(n833) );
  NAND20 U560 ( .A(n833), .B(n89), .Q(n12) );
  INV1 U561 ( .A(n683), .Q(n773) );
  XOR21 U562 ( .A(n30), .B(n785), .Q(SUM[8]) );
  CLKIN0 U563 ( .A(n98), .Q(n834) );
  NAND20 U564 ( .A(n171), .B(n815), .Q(n158) );
  NAND21 U565 ( .A(n841), .B(n62), .Q(n9) );
  NAND20 U566 ( .A(n823), .B(n231), .Q(n28) );
  NAND21 U567 ( .A(n815), .B(n163), .Q(n20) );
  INV3 U568 ( .A(n231), .Q(n822) );
  INV0 U569 ( .A(n126), .Q(n849) );
  NAND21 U570 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NOR20 U571 ( .A(n828), .B(n6), .Q(n55) );
  INV1 U572 ( .A(n6), .Q(n832) );
  AOI212 U573 ( .A(n764), .B(n179), .C(n180), .Q(n178) );
  AOI210 U574 ( .A(n775), .B(n825), .C(n204), .Q(n198) );
  INV2 U575 ( .A(n15), .Q(n809) );
  INV2 U576 ( .A(n21), .Q(n820) );
  NAND20 U577 ( .A(n798), .B(n771), .Q(n34) );
  CLKIN3 U578 ( .A(n59), .Q(n828) );
  INV0 U579 ( .A(n137), .Q(n812) );
  NAND20 U580 ( .A(n802), .B(n177), .Q(n22) );
  OAI210 U581 ( .A(n88), .B(n834), .C(n89), .Q(n85) );
  NAND20 U582 ( .A(n782), .B(n245), .Q(n30) );
  INV0 U583 ( .A(n61), .Q(n841) );
  INV0 U584 ( .A(n99), .Q(n835) );
  NAND21 U585 ( .A(n835), .B(n100), .Q(n13) );
  NAND20 U586 ( .A(n839), .B(n145), .Q(n18) );
  INV0 U587 ( .A(n255), .Q(n808) );
  INV0 U588 ( .A(n274), .Q(n789) );
  NAND20 U589 ( .A(n817), .B(n279), .Q(n37) );
  NAND20 U590 ( .A(n59), .B(n846), .Q(n46) );
  NAND20 U591 ( .A(n786), .B(n253), .Q(n31) );
  INV0 U592 ( .A(n117), .Q(n810) );
  INV3 U593 ( .A(n212), .Q(n843) );
  NAND21 U594 ( .A(B[14]), .B(A[14]), .Q(n195) );
  NAND20 U595 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U596 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U597 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV3 U598 ( .A(n53), .Q(n806) );
  INV3 U599 ( .A(n214), .Q(n776) );
  AOI211 U600 ( .A(n770), .B(n55), .C(n56), .Q(n769) );
  INV3 U601 ( .A(n60), .Q(n829) );
  INV3 U602 ( .A(n19), .Q(n818) );
  INV3 U603 ( .A(n16), .Q(n848) );
  NAND22 U604 ( .A(n842), .B(n776), .Q(n675) );
  INV3 U605 ( .A(n26), .Q(n842) );
  INV3 U606 ( .A(n29), .Q(n795) );
  NAND22 U607 ( .A(n804), .B(n839), .Q(n140) );
  INV3 U608 ( .A(n135), .Q(n813) );
  INV3 U609 ( .A(n171), .Q(n803) );
  INV3 U610 ( .A(n239), .Q(n783) );
  INV3 U611 ( .A(n771), .Q(n797) );
  INV3 U612 ( .A(n176), .Q(n802) );
  NAND20 U613 ( .A(n808), .B(n256), .Q(n32) );
  NAND20 U614 ( .A(n793), .B(n261), .Q(n33) );
  XOR21 U615 ( .A(n36), .B(n791), .Q(SUM[2]) );
  NAND20 U616 ( .A(n789), .B(n275), .Q(n36) );
  AOI210 U617 ( .A(n60), .B(n846), .C(n845), .Q(n47) );
  INV3 U618 ( .A(n51), .Q(n845) );
  NAND20 U619 ( .A(n138), .B(n812), .Q(n17) );
  NAND20 U620 ( .A(n826), .B(n206), .Q(n25) );
  NAND22 U621 ( .A(n784), .B(n843), .Q(n208) );
  NAND22 U622 ( .A(n807), .B(n195), .Q(n24) );
  NAND20 U623 ( .A(n794), .B(n186), .Q(n23) );
  INV0 U624 ( .A(n185), .Q(n794) );
  NAND22 U625 ( .A(n827), .B(n71), .Q(n10) );
  INV3 U626 ( .A(n70), .Q(n827) );
  INV0 U627 ( .A(n172), .Q(n799) );
  NAND22 U628 ( .A(n846), .B(n51), .Q(n8) );
  NAND22 U629 ( .A(n682), .B(n769), .Q(n52) );
  AOI210 U630 ( .A(n172), .B(n815), .C(n814), .Q(n159) );
  INV3 U631 ( .A(n163), .Q(n814) );
  NAND22 U632 ( .A(n830), .B(n80), .Q(n11) );
  INV3 U633 ( .A(n79), .Q(n830) );
  NOR21 U634 ( .A(n61), .B(n70), .Q(n59) );
  NAND22 U635 ( .A(n837), .B(n107), .Q(n14) );
  XOR21 U636 ( .A(n281), .B(n37), .Q(SUM[1]) );
  INV2 U637 ( .A(n278), .Q(n817) );
  NOR21 U638 ( .A(n70), .B(n6), .Q(n66) );
  NAND20 U639 ( .A(n821), .B(n174), .Q(n21) );
  INV3 U640 ( .A(n107), .Q(n838) );
  NAND21 U641 ( .A(n796), .B(n242), .Q(n29) );
  INV0 U642 ( .A(n241), .Q(n796) );
  NAND22 U643 ( .A(n849), .B(n127), .Q(n16) );
  NAND20 U644 ( .A(n810), .B(n118), .Q(n15) );
  NAND22 U645 ( .A(n819), .B(n156), .Q(n19) );
  AOI211 U646 ( .A(n775), .B(n843), .C(n844), .Q(n209) );
  INV3 U647 ( .A(n213), .Q(n844) );
  AOI211 U648 ( .A(n800), .B(n839), .C(n840), .Q(n141) );
  INV3 U649 ( .A(n145), .Q(n840) );
  NAND22 U650 ( .A(n500), .B(n21), .Q(n431) );
  INV3 U651 ( .A(n162), .Q(n815) );
  INV3 U652 ( .A(n144), .Q(n839) );
  BUF2 U653 ( .A(n266), .Q(n771) );
  NOR21 U654 ( .A(n88), .B(n836), .Q(n84) );
  NAND22 U655 ( .A(B[10]), .B(A[10]), .Q(n231) );
  NOR22 U656 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NAND22 U657 ( .A(A[16]), .B(B[16]), .Q(n177) );
  XNR21 U658 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U659 ( .A(n847), .B(n40), .Q(n7) );
  NAND22 U660 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR21 U661 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR22 U662 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND21 U663 ( .A(A[7]), .B(B[7]), .Q(n253) );
  INV3 U664 ( .A(n38), .Q(SUM[0]) );
  NAND22 U665 ( .A(n792), .B(n281), .Q(n38) );
  INV3 U666 ( .A(n280), .Q(n792) );
  NAND22 U667 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U668 ( .A(n50), .Q(n846) );
  NOR21 U669 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U670 ( .A(n39), .Q(n847) );
  NOR21 U671 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND21 U672 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND22 U673 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND21 U674 ( .A(n816), .B(n224), .Q(n27) );
  INV2 U675 ( .A(n194), .Q(n807) );
  OAI211 U676 ( .A(n194), .B(n824), .C(n195), .Q(n191) );
  NAND22 U678 ( .A(B[13]), .B(A[13]), .Q(n206) );
  NAND22 U679 ( .A(n119), .B(n15), .Q(n591) );
  NOR22 U680 ( .A(A[10]), .B(B[10]), .Q(n230) );
  NAND22 U681 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NOR22 U682 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR22 U683 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NAND22 U684 ( .A(B[9]), .B(A[9]), .Q(n242) );
  AOI210 U685 ( .A(n761), .B(n44), .C(n45), .Q(n43) );
endmodule


module adder_18 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_18_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_17_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n52, n53, n54, n57, n58, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n73, n74, n79, n80, n81, n82, n83, n84, n85, n88,
         n89, n90, n93, n94, n99, n100, n101, n102, n103, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n117, n118, n121,
         n122, n123, n124, n125, n126, n131, n132, n133, n134, n135, n139,
         n140, n141, n142, n147, n148, n149, n150, n151, n152, n153, n156,
         n157, n158, n161, n162, n167, n168, n169, n170, n171, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n186, n187, n188,
         n189, n194, n195, n196, n199, n200, n202, n203, n204, n205, n206,
         n207, n208, n209, n212, n213, n214, n215, n216, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n240, n241, n243, n244, n245, n246, n247, n248, n249,
         n250, n252, n253, n254, n255, n256, n391, n392, n393, n397, n398,
         n399, n400, n468, n469, n470, n475, n476, n545, n546, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830;

  OAI212 U16 ( .A(n53), .B(n45), .C(n46), .Q(n44) );
  OAI212 U32 ( .A(n770), .B(n761), .C(n769), .Q(n54) );
  OAI212 U36 ( .A(n771), .B(n74), .C(n772), .Q(n58) );
  OAI212 U46 ( .A(n66), .B(n761), .C(n67), .Q(n65) );
  OAI212 U70 ( .A(n84), .B(n761), .C(n85), .Q(n83) );
  OAI212 U80 ( .A(n785), .B(n761), .C(n786), .Q(n90) );
  OAI212 U242 ( .A(n208), .B(n817), .C(n209), .Q(n207) );
  OAI212 U252 ( .A(n215), .B(n817), .C(n216), .Q(n214) );
  OAI212 U263 ( .A(n223), .B(n243), .C(n224), .Q(n222) );
  OAI212 U267 ( .A(n231), .B(n227), .C(n228), .Q(n226) );
  OAI212 U273 ( .A(n230), .B(n232), .C(n231), .Q(n229) );
  OAI212 U281 ( .A(n241), .B(n235), .C(n236), .Q(n234) );
  OAI212 U298 ( .A(n250), .B(n246), .C(n247), .Q(n245) );
  OAI212 U304 ( .A(n249), .B(n815), .C(n250), .Q(n248) );
  OAI212 U311 ( .A(n256), .B(n253), .C(n254), .Q(n252) );
  OAI212 U324 ( .A(n174), .B(n202), .C(n175), .Q(n391) );
  OAI212 U337 ( .A(n759), .B(n795), .C(n171), .Q(n169) );
  OAI212 U373 ( .A(n810), .B(n795), .C(n808), .Q(n158) );
  OAI212 U368 ( .A(n152), .B(n795), .C(n153), .Q(n151) );
  OAI212 U355 ( .A(n186), .B(n178), .C(n179), .Q(n177) );
  OAI212 U384 ( .A(n107), .B(n142), .C(n108), .Q(n106) );
  AOI212 U401 ( .A(n391), .B(n105), .C(n106), .Q(n1) );
  AOI212 U376 ( .A(n147), .B(n397), .C(n148), .Q(n393) );
  OAI212 U396 ( .A(n71), .B(n63), .C(n64), .Q(n62) );
  OAI212 U435 ( .A(n171), .B(n167), .C(n168), .Q(n397) );
  OAI212 U378 ( .A(n114), .B(n795), .C(n115), .Q(n113) );
  AOI212 U432 ( .A(n189), .B(n176), .C(n177), .Q(n175) );
  OAI212 U367 ( .A(n765), .B(n761), .C(n764), .Q(n36) );
  OAI212 U365 ( .A(n183), .B(n797), .C(n760), .Q(n182) );
  OAI212 U420 ( .A(n209), .B(n205), .C(n206), .Q(n204) );
  OAI212 U441 ( .A(n48), .B(n761), .C(n49), .Q(n47) );
  NOR22 U325 ( .A(B[18]), .B(A[18]), .Q(n149) );
  NAND22 U326 ( .A(A[12]), .B(B[12]), .Q(n195) );
  INV0 U327 ( .A(n205), .Q(n806) );
  NOR24 U328 ( .A(B[10]), .B(A[10]), .Q(n205) );
  NOR22 U329 ( .A(n208), .B(n205), .Q(n203) );
  AOI212 U330 ( .A(n807), .B(n188), .C(n189), .Q(n187) );
  CLKIN6 U331 ( .A(n202), .Q(n807) );
  XOR22 U332 ( .A(n187), .B(n20), .Q(SUM[13]) );
  NOR24 U333 ( .A(B[20]), .B(A[20]), .Q(n131) );
  NAND22 U334 ( .A(A[19]), .B(B[19]), .Q(n139) );
  NOR23 U335 ( .A(n771), .B(n73), .Q(n57) );
  XNR22 U336 ( .A(n17), .B(n169), .Q(SUM[16]) );
  XNR22 U338 ( .A(n9), .B(n101), .Q(SUM[24]) );
  XNR22 U339 ( .A(n15), .B(n151), .Q(SUM[18]) );
  XOR22 U340 ( .A(n18), .B(n795), .Q(SUM[15]) );
  NAND26 U341 ( .A(A[11]), .B(B[11]), .Q(n200) );
  NOR23 U342 ( .A(B[11]), .B(A[11]), .Q(n199) );
  NOR21 U343 ( .A(B[15]), .B(A[15]), .Q(n170) );
  NAND24 U344 ( .A(n147), .B(n161), .Q(n141) );
  INV1 U345 ( .A(n156), .Q(n813) );
  NAND24 U346 ( .A(A[15]), .B(B[15]), .Q(n171) );
  NOR21 U347 ( .A(B[15]), .B(A[15]), .Q(n759) );
  NAND23 U348 ( .A(A[16]), .B(B[16]), .Q(n168) );
  NAND23 U349 ( .A(n470), .B(n150), .Q(n148) );
  NOR22 U350 ( .A(n149), .B(n156), .Q(n147) );
  INV3 U351 ( .A(n73), .Q(n776) );
  NOR23 U352 ( .A(B[21]), .B(A[21]), .Q(n118) );
  NOR21 U353 ( .A(n99), .B(n102), .Q(n93) );
  NAND22 U354 ( .A(n93), .B(n79), .Q(n73) );
  NAND22 U356 ( .A(A[20]), .B(B[20]), .Q(n132) );
  INV3 U357 ( .A(n118), .Q(n802) );
  NAND24 U358 ( .A(n545), .B(n546), .Q(SUM[19]) );
  CLKIN3 U359 ( .A(n178), .Q(n799) );
  NAND22 U360 ( .A(n802), .B(n125), .Q(n392) );
  OAI211 U361 ( .A(n141), .B(n795), .C(n393), .Q(n140) );
  NAND23 U362 ( .A(n780), .B(n803), .Q(n546) );
  NAND20 U363 ( .A(n804), .B(n139), .Q(n14) );
  INV3 U364 ( .A(n400), .Q(n804) );
  NAND21 U366 ( .A(A[13]), .B(B[13]), .Q(n186) );
  NOR21 U369 ( .A(B[30]), .B(A[30]), .Q(n45) );
  AOI212 U370 ( .A(n162), .B(n147), .C(n148), .Q(n142) );
  CLKIN0 U371 ( .A(n139), .Q(n805) );
  OAI211 U372 ( .A(n139), .B(n131), .C(n132), .Q(n126) );
  OAI211 U374 ( .A(n139), .B(n131), .C(n132), .Q(n399) );
  XNR22 U375 ( .A(n4), .B(n54), .Q(SUM[29]) );
  XNR22 U377 ( .A(n3), .B(n47), .Q(SUM[30]) );
  NOR24 U379 ( .A(B[13]), .B(A[13]), .Q(n183) );
  XNR22 U380 ( .A(n13), .B(n133), .Q(SUM[20]) );
  OAI211 U381 ( .A(n134), .B(n795), .C(n135), .Q(n133) );
  XNR22 U382 ( .A(n5), .B(n65), .Q(SUM[28]) );
  AOI212 U383 ( .A(n126), .B(n109), .C(n110), .Q(n108) );
  OAI212 U385 ( .A(n121), .B(n111), .C(n112), .Q(n110) );
  NAND21 U386 ( .A(A[22]), .B(B[22]), .Q(n112) );
  NOR22 U387 ( .A(B[19]), .B(A[19]), .Q(n400) );
  AOI212 U388 ( .A(n807), .B(n181), .C(n182), .Q(n180) );
  NOR21 U389 ( .A(n183), .B(n794), .Q(n181) );
  XNR22 U390 ( .A(n16), .B(n158), .Q(SUM[17]) );
  CLKIN4 U391 ( .A(n149), .Q(n781) );
  XNR22 U392 ( .A(n12), .B(n122), .Q(SUM[21]) );
  XNR22 U393 ( .A(n6), .B(n72), .Q(SUM[27]) );
  XOR22 U394 ( .A(n19), .B(n180), .Q(SUM[14]) );
  NOR21 U395 ( .A(B[28]), .B(A[28]), .Q(n63) );
  NAND22 U397 ( .A(n787), .B(n89), .Q(n8) );
  NAND21 U398 ( .A(A[25]), .B(B[25]), .Q(n89) );
  NOR22 U399 ( .A(n81), .B(n88), .Q(n79) );
  NOR21 U400 ( .A(B[25]), .B(A[25]), .Q(n88) );
  OAI211 U402 ( .A(n89), .B(n81), .C(n82), .Q(n80) );
  NOR24 U403 ( .A(B[22]), .B(A[22]), .Q(n111) );
  NAND21 U404 ( .A(n783), .B(n761), .Q(n476) );
  BUF15 U405 ( .A(n1), .Q(n761) );
  NAND21 U406 ( .A(A[18]), .B(B[18]), .Q(n150) );
  XNR22 U407 ( .A(n7), .B(n83), .Q(SUM[26]) );
  NAND21 U408 ( .A(A[14]), .B(B[14]), .Q(n179) );
  OAI212 U409 ( .A(n200), .B(n194), .C(n195), .Q(n189) );
  NOR24 U410 ( .A(B[12]), .B(A[12]), .Q(n194) );
  CLKIN2 U411 ( .A(n189), .Q(n797) );
  AOI212 U412 ( .A(n94), .B(n79), .C(n80), .Q(n74) );
  NOR24 U413 ( .A(B[17]), .B(A[17]), .Q(n156) );
  XNR22 U414 ( .A(n11), .B(n113), .Q(SUM[22]) );
  NOR21 U415 ( .A(B[26]), .B(A[26]), .Q(n81) );
  OAI212 U416 ( .A(n73), .B(n761), .C(n74), .Q(n72) );
  NOR20 U417 ( .A(n41), .B(n73), .Q(n39) );
  OAI212 U418 ( .A(n103), .B(n99), .C(n100), .Q(n94) );
  OAI212 U419 ( .A(n102), .B(n761), .C(n103), .Q(n101) );
  NAND22 U421 ( .A(A[23]), .B(B[23]), .Q(n103) );
  OAI210 U422 ( .A(n41), .B(n74), .C(n42), .Q(n40) );
  NOR23 U423 ( .A(n167), .B(n170), .Q(n161) );
  INV1 U424 ( .A(n167), .Q(n811) );
  OAI211 U425 ( .A(n171), .B(n167), .C(n168), .Q(n398) );
  OAI211 U426 ( .A(n171), .B(n167), .C(n168), .Q(n162) );
  NOR24 U427 ( .A(B[16]), .B(A[16]), .Q(n167) );
  NOR22 U428 ( .A(n111), .B(n118), .Q(n109) );
  NAND22 U429 ( .A(A[17]), .B(B[17]), .Q(n157) );
  OAI211 U430 ( .A(n118), .B(n791), .C(n121), .Q(n117) );
  NAND22 U431 ( .A(n802), .B(n121), .Q(n12) );
  NAND21 U433 ( .A(A[21]), .B(B[21]), .Q(n121) );
  INV1 U434 ( .A(n81), .Q(n775) );
  NOR22 U436 ( .A(B[23]), .B(A[23]), .Q(n102) );
  NOR23 U437 ( .A(n131), .B(n400), .Q(n125) );
  XNR22 U438 ( .A(n8), .B(n90), .Q(SUM[25]) );
  NOR21 U439 ( .A(B[24]), .B(A[24]), .Q(n99) );
  OAI211 U440 ( .A(n123), .B(n795), .C(n124), .Q(n122) );
  NAND21 U442 ( .A(n782), .B(n125), .Q(n123) );
  NAND20 U443 ( .A(A[13]), .B(B[13]), .Q(n760) );
  INV3 U444 ( .A(n759), .Q(n809) );
  INV3 U445 ( .A(n393), .Q(n779) );
  NAND22 U446 ( .A(n475), .B(n476), .Q(SUM[23]) );
  NAND20 U447 ( .A(n93), .B(n787), .Q(n84) );
  NOR22 U448 ( .A(n107), .B(n141), .Q(n105) );
  CLKIN3 U449 ( .A(n58), .Q(n769) );
  INV2 U450 ( .A(n74), .Q(n777) );
  CLKIN3 U451 ( .A(n40), .Q(n764) );
  INV0 U452 ( .A(n45), .Q(n763) );
  NOR22 U453 ( .A(B[14]), .B(A[14]), .Q(n178) );
  NAND21 U454 ( .A(n57), .B(n767), .Q(n48) );
  NAND22 U455 ( .A(n10), .B(n778), .Q(n475) );
  NAND22 U456 ( .A(n768), .B(n64), .Q(n5) );
  INV0 U457 ( .A(n63), .Q(n768) );
  INV2 U458 ( .A(n399), .Q(n791) );
  AOI210 U459 ( .A(n779), .B(n792), .C(n117), .Q(n115) );
  INV2 U460 ( .A(n469), .Q(n773) );
  NAND20 U461 ( .A(n798), .B(n112), .Q(n11) );
  CLKIN0 U462 ( .A(n93), .Q(n785) );
  NOR21 U463 ( .A(n45), .B(n52), .Q(n43) );
  XNR21 U464 ( .A(n22), .B(n807), .Q(SUM[11]) );
  NAND20 U465 ( .A(A[4]), .B(B[4]), .Q(n241) );
  NAND20 U466 ( .A(A[8]), .B(B[8]), .Q(n216) );
  NAND20 U467 ( .A(A[9]), .B(B[9]), .Q(n213) );
  NAND21 U468 ( .A(n782), .B(n792), .Q(n114) );
  AOI210 U469 ( .A(n779), .B(n125), .C(n399), .Q(n124) );
  NAND20 U470 ( .A(n161), .B(n813), .Q(n152) );
  NAND20 U471 ( .A(n61), .B(n43), .Q(n41) );
  NOR22 U472 ( .A(n194), .B(n199), .Q(n188) );
  NAND20 U473 ( .A(n809), .B(n171), .Q(n18) );
  NOR22 U474 ( .A(n183), .B(n178), .Q(n176) );
  INV0 U475 ( .A(n183), .Q(n801) );
  CLKIN0 U476 ( .A(n161), .Q(n810) );
  INV0 U477 ( .A(n111), .Q(n798) );
  AOI210 U478 ( .A(n398), .B(n813), .C(n812), .Q(n153) );
  NAND20 U479 ( .A(n150), .B(n781), .Q(n15) );
  AOI212 U480 ( .A(n203), .B(n222), .C(n204), .Q(n202) );
  NAND20 U481 ( .A(n806), .B(n206), .Q(n23) );
  AOI210 U482 ( .A(n62), .B(n43), .C(n44), .Q(n42) );
  INV0 U483 ( .A(n199), .Q(n793) );
  AOI211 U484 ( .A(n779), .B(n804), .C(n805), .Q(n135) );
  NAND20 U485 ( .A(A[29]), .B(B[29]), .Q(n53) );
  NAND20 U486 ( .A(A[27]), .B(B[27]), .Q(n469) );
  NAND20 U487 ( .A(A[26]), .B(B[26]), .Q(n82) );
  NOR20 U488 ( .A(B[27]), .B(A[27]), .Q(n70) );
  INV3 U489 ( .A(n140), .Q(n780) );
  INV3 U490 ( .A(n141), .Q(n782) );
  INV3 U491 ( .A(n761), .Q(n778) );
  INV3 U492 ( .A(n39), .Q(n765) );
  INV6 U493 ( .A(n391), .Q(n795) );
  NAND22 U494 ( .A(n140), .B(n14), .Q(n545) );
  INV3 U495 ( .A(n14), .Q(n803) );
  INV3 U496 ( .A(n10), .Q(n783) );
  NAND22 U497 ( .A(n125), .B(n109), .Q(n107) );
  NAND22 U498 ( .A(n776), .B(n774), .Q(n66) );
  NAND22 U499 ( .A(n782), .B(n804), .Q(n134) );
  INV3 U500 ( .A(n392), .Q(n792) );
  INV3 U501 ( .A(n61), .Q(n771) );
  INV0 U502 ( .A(n397), .Q(n808) );
  AOI211 U503 ( .A(n816), .B(n233), .C(n234), .Q(n232) );
  INV3 U504 ( .A(n222), .Q(n817) );
  INV3 U505 ( .A(n243), .Q(n816) );
  INV3 U506 ( .A(n252), .Q(n815) );
  XOR21 U507 ( .A(n21), .B(n196), .Q(SUM[12]) );
  NAND22 U508 ( .A(n800), .B(n195), .Q(n21) );
  AOI211 U509 ( .A(n807), .B(n793), .C(n796), .Q(n196) );
  INV3 U510 ( .A(n194), .Q(n800) );
  NAND22 U511 ( .A(n799), .B(n179), .Q(n19) );
  NAND22 U512 ( .A(n790), .B(n132), .Q(n13) );
  INV3 U513 ( .A(n131), .Q(n790) );
  NAND22 U514 ( .A(n767), .B(n53), .Q(n4) );
  CLKIN3 U515 ( .A(n57), .Q(n770) );
  NAND22 U516 ( .A(n793), .B(n200), .Q(n22) );
  XNR21 U517 ( .A(n23), .B(n207), .Q(SUM[10]) );
  INV3 U518 ( .A(n62), .Q(n772) );
  NAND22 U519 ( .A(n188), .B(n176), .Q(n174) );
  NAND22 U520 ( .A(n763), .B(n46), .Q(n3) );
  NAND22 U521 ( .A(n811), .B(n168), .Q(n17) );
  NAND22 U522 ( .A(n775), .B(n82), .Q(n7) );
  NAND22 U523 ( .A(n774), .B(n469), .Q(n6) );
  NOR21 U524 ( .A(n63), .B(n70), .Q(n61) );
  NAND22 U525 ( .A(n813), .B(n157), .Q(n16) );
  NAND22 U526 ( .A(n801), .B(n760), .Q(n20) );
  AOI210 U527 ( .A(n94), .B(n787), .C(n788), .Q(n85) );
  INV3 U528 ( .A(n89), .Q(n788) );
  NAND22 U529 ( .A(n784), .B(n103), .Q(n10) );
  INV3 U530 ( .A(n102), .Q(n784) );
  AOI210 U531 ( .A(n58), .B(n767), .C(n766), .Q(n49) );
  INV3 U532 ( .A(n53), .Q(n766) );
  NAND22 U533 ( .A(n812), .B(n781), .Q(n470) );
  INV3 U534 ( .A(n70), .Q(n774) );
  INV3 U535 ( .A(n88), .Q(n787) );
  INV3 U536 ( .A(n52), .Q(n767) );
  AOI211 U537 ( .A(n777), .B(n774), .C(n773), .Q(n67) );
  INV0 U538 ( .A(n94), .Q(n786) );
  INV3 U539 ( .A(n157), .Q(n812) );
  INV3 U540 ( .A(n99), .Q(n789) );
  CLKIN0 U541 ( .A(n188), .Q(n794) );
  INV3 U542 ( .A(n200), .Q(n796) );
  XOR21 U543 ( .A(n28), .B(n237), .Q(SUM[5]) );
  NAND22 U544 ( .A(n824), .B(n236), .Q(n28) );
  AOI211 U545 ( .A(n816), .B(n823), .C(n822), .Q(n237) );
  INV3 U546 ( .A(n235), .Q(n824) );
  XOR21 U547 ( .A(n31), .B(n815), .Q(SUM[2]) );
  NAND22 U548 ( .A(n820), .B(n250), .Q(n31) );
  INV3 U549 ( .A(n249), .Q(n820) );
  XOR21 U550 ( .A(n27), .B(n232), .Q(SUM[6]) );
  NAND22 U551 ( .A(n825), .B(n231), .Q(n27) );
  INV3 U552 ( .A(n230), .Q(n825) );
  XOR21 U553 ( .A(n25), .B(n817), .Q(SUM[8]) );
  NAND22 U554 ( .A(n828), .B(n216), .Q(n25) );
  NAND22 U555 ( .A(n233), .B(n225), .Q(n223) );
  AOI211 U556 ( .A(n234), .B(n225), .C(n226), .Q(n224) );
  NOR21 U557 ( .A(n227), .B(n230), .Q(n225) );
  AOI211 U558 ( .A(n252), .B(n244), .C(n245), .Q(n243) );
  NOR21 U559 ( .A(n246), .B(n249), .Q(n244) );
  XNR21 U560 ( .A(n24), .B(n214), .Q(SUM[9]) );
  NAND22 U561 ( .A(n830), .B(n213), .Q(n24) );
  XNR21 U562 ( .A(n29), .B(n816), .Q(SUM[4]) );
  NAND22 U563 ( .A(n823), .B(n241), .Q(n29) );
  XNR21 U564 ( .A(n26), .B(n229), .Q(SUM[7]) );
  NAND22 U565 ( .A(n826), .B(n228), .Q(n26) );
  INV3 U566 ( .A(n227), .Q(n826) );
  XNR21 U567 ( .A(n30), .B(n248), .Q(SUM[3]) );
  NAND22 U568 ( .A(n821), .B(n247), .Q(n30) );
  INV3 U569 ( .A(n246), .Q(n821) );
  XOR21 U570 ( .A(n256), .B(n32), .Q(SUM[1]) );
  NAND22 U571 ( .A(n819), .B(n254), .Q(n32) );
  INV3 U572 ( .A(n253), .Q(n819) );
  AOI211 U573 ( .A(n830), .B(n827), .C(n829), .Q(n209) );
  INV3 U574 ( .A(n213), .Q(n829) );
  INV3 U575 ( .A(n216), .Q(n827) );
  NOR21 U576 ( .A(n235), .B(n240), .Q(n233) );
  NAND22 U577 ( .A(n828), .B(n830), .Q(n208) );
  INV3 U578 ( .A(n215), .Q(n828) );
  INV3 U579 ( .A(n240), .Q(n823) );
  INV3 U580 ( .A(n241), .Q(n822) );
  NAND20 U581 ( .A(A[24]), .B(B[24]), .Q(n100) );
  NAND22 U582 ( .A(n789), .B(n468), .Q(n9) );
  NAND20 U583 ( .A(A[24]), .B(B[24]), .Q(n468) );
  XNR21 U584 ( .A(n2), .B(n36), .Q(SUM[31]) );
  NAND22 U585 ( .A(n762), .B(n35), .Q(n2) );
  NAND20 U586 ( .A(A[31]), .B(B[31]), .Q(n35) );
  NAND20 U587 ( .A(A[27]), .B(B[27]), .Q(n71) );
  NOR20 U588 ( .A(B[29]), .B(A[29]), .Q(n52) );
  NAND22 U589 ( .A(A[10]), .B(B[10]), .Q(n206) );
  NAND20 U590 ( .A(A[28]), .B(B[28]), .Q(n64) );
  INV3 U591 ( .A(n34), .Q(n762) );
  NOR20 U592 ( .A(B[31]), .B(A[31]), .Q(n34) );
  NAND20 U593 ( .A(A[30]), .B(B[30]), .Q(n46) );
  NOR20 U594 ( .A(B[7]), .B(A[7]), .Q(n227) );
  NOR20 U595 ( .A(B[5]), .B(A[5]), .Q(n235) );
  NOR20 U596 ( .A(B[3]), .B(A[3]), .Q(n246) );
  NOR20 U597 ( .A(B[6]), .B(A[6]), .Q(n230) );
  NOR20 U598 ( .A(B[2]), .B(A[2]), .Q(n249) );
  NOR20 U599 ( .A(B[4]), .B(A[4]), .Q(n240) );
  NOR20 U600 ( .A(B[1]), .B(A[1]), .Q(n253) );
  NOR20 U601 ( .A(B[8]), .B(A[8]), .Q(n215) );
  NAND20 U602 ( .A(A[0]), .B(B[0]), .Q(n256) );
  NAND20 U603 ( .A(A[6]), .B(B[6]), .Q(n231) );
  NAND20 U604 ( .A(A[2]), .B(B[2]), .Q(n250) );
  NAND20 U605 ( .A(A[1]), .B(B[1]), .Q(n254) );
  NAND20 U606 ( .A(A[7]), .B(B[7]), .Q(n228) );
  NAND20 U607 ( .A(A[5]), .B(B[5]), .Q(n236) );
  NAND20 U608 ( .A(A[3]), .B(B[3]), .Q(n247) );
  INV3 U609 ( .A(n212), .Q(n830) );
  NOR20 U610 ( .A(B[9]), .B(A[9]), .Q(n212) );
  INV3 U611 ( .A(n33), .Q(SUM[0]) );
  NAND22 U612 ( .A(n818), .B(n256), .Q(n33) );
  INV3 U613 ( .A(n255), .Q(n818) );
  NOR20 U614 ( .A(B[0]), .B(A[0]), .Q(n255) );
endmodule


module adder_17 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_17_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module reg_5 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30,
         n32, n35, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n53, n54, n55, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n104, n105, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393;

  DF3 Dout_reg_16_ ( .D(n71), .C(Clk), .Q(Dout[16]), .QN(n4) );
  DF3 Dout_reg_15_ ( .D(n85), .C(Clk), .Q(Dout[15]), .QN(n73) );
  DF3 Dout_reg_14_ ( .D(n86), .C(Clk), .Q(Dout[14]), .QN(n72) );
  DF3 Dout_reg_13_ ( .D(n87), .C(Clk), .Q(Dout[13]), .QN(n55) );
  DF3 Dout_reg_12_ ( .D(n88), .C(Clk), .Q(Dout[12]), .QN(n53) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n77) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n75) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n74) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n81) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n80) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n79) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n78) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n84) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n83) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n82) );
  DF3 Dout_reg_11_ ( .D(n89), .C(Clk), .Q(Dout[11]), .QN(n54) );
  DF3 Dout_reg_23_ ( .D(n64), .C(Clk), .Q(Dout[23]), .QN(n18) );
  DF3 Dout_reg_25_ ( .D(n62), .C(Clk), .Q(Dout[25]), .QN(n22) );
  DF3 Dout_reg_22_ ( .D(n65), .C(Clk), .Q(Dout[22]), .QN(n16) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n76) );
  OAI222 U3 ( .A(n83), .B(n358), .C(n360), .D(n392), .Q(n99) );
  OAI222 U4 ( .A(n84), .B(n358), .C(n359), .D(n393), .Q(n98) );
  OAI222 U5 ( .A(n78), .B(n358), .C(n104), .D(n388), .Q(n97) );
  OAI222 U6 ( .A(n79), .B(n358), .C(n360), .D(n390), .Q(n96) );
  OAI222 U7 ( .A(n80), .B(n358), .C(n359), .D(n389), .Q(n95) );
  OAI222 U8 ( .A(n81), .B(n358), .C(n104), .D(n387), .Q(n94) );
  OAI222 U9 ( .A(n74), .B(n358), .C(n360), .D(n386), .Q(n93) );
  OAI222 U10 ( .A(n75), .B(n358), .C(n359), .D(n384), .Q(n92) );
  OAI222 U11 ( .A(n76), .B(n358), .C(n104), .D(n385), .Q(n91) );
  OAI222 U12 ( .A(n77), .B(n358), .C(n360), .D(n383), .Q(n90) );
  OAI222 U13 ( .A(n54), .B(n358), .C(n359), .D(n382), .Q(n89) );
  OAI222 U14 ( .A(n53), .B(n358), .C(n104), .D(n381), .Q(n88) );
  OAI222 U15 ( .A(n55), .B(n358), .C(n360), .D(n379), .Q(n87) );
  OAI222 U16 ( .A(n72), .B(n358), .C(n359), .D(n380), .Q(n86) );
  OAI222 U17 ( .A(n73), .B(n358), .C(n104), .D(n376), .Q(n85) );
  OAI222 U18 ( .A(n4), .B(n358), .C(n360), .D(n378), .Q(n71) );
  OAI222 U19 ( .A(n6), .B(n358), .C(n377), .D(n359), .Q(n70) );
  OAI222 U20 ( .A(n8), .B(n358), .C(n104), .D(n375), .Q(n69) );
  OAI222 U21 ( .A(n10), .B(n358), .C(n360), .D(n370), .Q(n68) );
  OAI222 U22 ( .A(n12), .B(n358), .C(n359), .D(n374), .Q(n67) );
  OAI222 U23 ( .A(n14), .B(n358), .C(n104), .D(n371), .Q(n66) );
  OAI222 U24 ( .A(n16), .B(n358), .C(n360), .D(n373), .Q(n65) );
  OAI222 U25 ( .A(n18), .B(n358), .C(n372), .D(n359), .Q(n64) );
  OAI222 U26 ( .A(n20), .B(n358), .C(n104), .D(n369), .Q(n63) );
  OAI222 U27 ( .A(n22), .B(n358), .C(n360), .D(n368), .Q(n62) );
  OAI222 U28 ( .A(n24), .B(n358), .C(n359), .D(n367), .Q(n61) );
  OAI222 U29 ( .A(n26), .B(n358), .C(n104), .D(n366), .Q(n60) );
  OAI222 U30 ( .A(n28), .B(n358), .C(n360), .D(n365), .Q(n59) );
  OAI222 U31 ( .A(n30), .B(n358), .C(n359), .D(n364), .Q(n58) );
  OAI222 U32 ( .A(n32), .B(n358), .C(n104), .D(n363), .Q(n57) );
  OAI222 U33 ( .A(n35), .B(n358), .C(n360), .D(n362), .Q(n56) );
  OAI222 U34 ( .A(n82), .B(n358), .C(n359), .D(n391), .Q(n100) );
  DF1 Dout_reg_30_ ( .D(n57), .C(Clk), .Q(Dout[30]), .QN(n32) );
  DF1 Dout_reg_27_ ( .D(n60), .C(Clk), .Q(Dout[27]), .QN(n26) );
  DF1 Dout_reg_28_ ( .D(n59), .C(Clk), .Q(Dout[28]), .QN(n28) );
  DF1 Dout_reg_20_ ( .D(n67), .C(Clk), .Q(Dout[20]), .QN(n12) );
  DF1 Dout_reg_21_ ( .D(n66), .C(Clk), .Q(Dout[21]), .QN(n14) );
  DF1 Dout_reg_24_ ( .D(n63), .C(Clk), .Q(Dout[24]), .QN(n20) );
  DF1 Dout_reg_18_ ( .D(n69), .C(Clk), .Q(Dout[18]), .QN(n8) );
  DF1 Dout_reg_17_ ( .D(n70), .C(Clk), .Q(Dout[17]), .QN(n6) );
  DF1 Dout_reg_19_ ( .D(n68), .C(Clk), .Q(Dout[19]), .QN(n10) );
  DF1 Dout_reg_31_ ( .D(n56), .C(Clk), .Q(Dout[31]), .QN(n35) );
  DF1 Dout_reg_26_ ( .D(n61), .C(Clk), .Q(Dout[26]), .QN(n24) );
  DF3 Dout_reg_29_ ( .D(n58), .C(Clk), .Q(Dout[29]), .QN(n30) );
  INV3 U35 ( .A(Din[24]), .Q(n369) );
  INV4 U36 ( .A(Din[26]), .Q(n367) );
  INV4 U37 ( .A(Din[25]), .Q(n368) );
  INV3 U38 ( .A(Din[19]), .Q(n370) );
  INV3 U39 ( .A(Din[18]), .Q(n375) );
  INV3 U40 ( .A(Din[21]), .Q(n371) );
  INV3 U41 ( .A(Din[9]), .Q(n385) );
  INV4 U42 ( .A(Din[27]), .Q(n366) );
  INV3 U43 ( .A(Din[29]), .Q(n364) );
  INV3 U44 ( .A(Din[30]), .Q(n363) );
  INV3 U45 ( .A(Din[31]), .Q(n362) );
  INV3 U46 ( .A(Din[20]), .Q(n374) );
  INV4 U47 ( .A(Din[28]), .Q(n365) );
  INV3 U48 ( .A(Din[17]), .Q(n377) );
  INV3 U49 ( .A(Din[23]), .Q(n372) );
  INV3 U50 ( .A(Din[22]), .Q(n373) );
  INV2 U51 ( .A(Din[13]), .Q(n379) );
  INV2 U52 ( .A(Din[11]), .Q(n382) );
  INV2 U53 ( .A(Din[14]), .Q(n380) );
  CLKIN3 U54 ( .A(Din[8]), .Q(n384) );
  INV2 U55 ( .A(Din[10]), .Q(n383) );
  CLKIN3 U56 ( .A(Din[7]), .Q(n386) );
  INV2 U57 ( .A(Din[15]), .Q(n376) );
  NAND22 U58 ( .A(n361), .B(n358), .Q(n359) );
  NAND22 U59 ( .A(n361), .B(n358), .Q(n360) );
  NAND22 U60 ( .A(n361), .B(n358), .Q(n104) );
  INV3 U61 ( .A(Reset), .Q(n361) );
  INV3 U62 ( .A(n105), .Q(n358) );
  INV3 U63 ( .A(Din[12]), .Q(n381) );
  CLKIN3 U64 ( .A(Din[16]), .Q(n378) );
  INV3 U65 ( .A(Din[3]), .Q(n388) );
  INV3 U66 ( .A(Din[4]), .Q(n390) );
  INV3 U67 ( .A(Din[6]), .Q(n387) );
  INV3 U68 ( .A(Din[5]), .Q(n389) );
  INV3 U69 ( .A(Din[0]), .Q(n391) );
  INV3 U70 ( .A(Din[1]), .Q(n392) );
  INV3 U71 ( .A(Din[2]), .Q(n393) );
  NOR21 U72 ( .A(Load), .B(Reset), .Q(n105) );
endmodule


module reg_4 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32,
         n35, n47, n49, n51, n53, n55, n57, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n58, n59, n60, n61, n62, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n104, n105, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398;

  DF3 Dout_reg_16_ ( .D(n78), .C(Clk), .Q(Dout[16]), .QN(n16) );
  DF3 Dout_reg_15_ ( .D(n79), .C(Clk), .Q(Dout[15]), .QN(n14) );
  DF3 Dout_reg_14_ ( .D(n80), .C(Clk), .Q(Dout[14]), .QN(n12) );
  DF3 Dout_reg_12_ ( .D(n82), .C(Clk), .Q(Dout[12]), .QN(n8) );
  DF3 Dout_reg_11_ ( .D(n83), .C(Clk), .Q(Dout[11]), .QN(n6) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n58) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n59) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n85) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n62) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n61) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n87) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n86) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n84) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n89) );
  DF3 Dout_reg_13_ ( .D(n81), .C(Clk), .Q(Dout[13]), .QN(n10) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n88) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n60) );
  DF3 Dout_reg_21_ ( .D(n73), .C(Clk), .Q(Dout[21]), .QN(n26) );
  OAI222 U3 ( .A(n88), .B(n363), .C(n365), .D(n394), .Q(n99) );
  OAI222 U4 ( .A(n87), .B(n363), .C(n364), .D(n397), .Q(n98) );
  OAI222 U5 ( .A(n86), .B(n363), .C(n104), .D(n396), .Q(n97) );
  OAI222 U6 ( .A(n61), .B(n363), .C(n365), .D(n398), .Q(n96) );
  OAI222 U7 ( .A(n62), .B(n363), .C(n364), .D(n388), .Q(n95) );
  OAI222 U8 ( .A(n85), .B(n363), .C(n104), .D(n390), .Q(n94) );
  OAI222 U9 ( .A(n84), .B(n363), .C(n365), .D(n389), .Q(n93) );
  OAI222 U10 ( .A(n59), .B(n363), .C(n364), .D(n392), .Q(n92) );
  OAI222 U11 ( .A(n60), .B(n363), .C(n104), .D(n393), .Q(n91) );
  OAI222 U12 ( .A(n58), .B(n363), .C(n365), .D(n391), .Q(n90) );
  OAI222 U13 ( .A(n6), .B(n363), .C(n364), .D(n387), .Q(n83) );
  OAI222 U14 ( .A(n8), .B(n363), .C(n104), .D(n386), .Q(n82) );
  OAI222 U15 ( .A(n10), .B(n363), .C(n365), .D(n385), .Q(n81) );
  OAI222 U16 ( .A(n12), .B(n363), .C(n364), .D(n383), .Q(n80) );
  OAI222 U17 ( .A(n14), .B(n363), .C(n104), .D(n384), .Q(n79) );
  OAI222 U18 ( .A(n16), .B(n363), .C(n365), .D(n382), .Q(n78) );
  OAI222 U19 ( .A(n18), .B(n363), .C(n364), .D(n381), .Q(n77) );
  OAI222 U20 ( .A(n20), .B(n363), .C(n104), .D(n380), .Q(n76) );
  OAI222 U21 ( .A(n22), .B(n363), .C(n365), .D(n379), .Q(n75) );
  OAI222 U22 ( .A(n24), .B(n363), .C(n364), .D(n378), .Q(n74) );
  OAI222 U23 ( .A(n26), .B(n363), .C(n104), .D(n375), .Q(n73) );
  OAI222 U24 ( .A(n28), .B(n363), .C(n365), .D(n377), .Q(n72) );
  OAI222 U25 ( .A(n30), .B(n363), .C(n364), .D(n376), .Q(n71) );
  OAI222 U26 ( .A(n32), .B(n363), .C(n104), .D(n374), .Q(n70) );
  OAI222 U27 ( .A(n35), .B(n363), .C(n365), .D(n373), .Q(n69) );
  OAI222 U28 ( .A(n47), .B(n363), .C(n364), .D(n372), .Q(n68) );
  OAI222 U29 ( .A(n49), .B(n363), .C(n104), .D(n371), .Q(n67) );
  OAI222 U30 ( .A(n51), .B(n363), .C(n365), .D(n370), .Q(n66) );
  OAI222 U31 ( .A(n53), .B(n363), .C(n364), .D(n369), .Q(n65) );
  OAI222 U32 ( .A(n55), .B(n363), .C(n104), .D(n368), .Q(n64) );
  OAI222 U33 ( .A(n57), .B(n363), .C(n365), .D(n367), .Q(n63) );
  OAI222 U34 ( .A(n89), .B(n363), .C(n364), .D(n395), .Q(n100) );
  DF1 Dout_reg_27_ ( .D(n67), .C(Clk), .Q(Dout[27]), .QN(n49) );
  DF1 Dout_reg_30_ ( .D(n64), .C(Clk), .Q(Dout[30]), .QN(n55) );
  DF1 Dout_reg_23_ ( .D(n71), .C(Clk), .Q(Dout[23]), .QN(n30) );
  DF1 Dout_reg_22_ ( .D(n72), .C(Clk), .Q(Dout[22]), .QN(n28) );
  DF1 Dout_reg_18_ ( .D(n76), .C(Clk), .Q(Dout[18]), .QN(n20) );
  DF1 Dout_reg_29_ ( .D(n65), .C(Clk), .Q(Dout[29]), .QN(n53) );
  DF1 Dout_reg_20_ ( .D(n74), .C(Clk), .Q(Dout[20]), .QN(n24) );
  DF1 Dout_reg_19_ ( .D(n75), .C(Clk), .Q(Dout[19]), .QN(n22) );
  DF1 Dout_reg_24_ ( .D(n70), .C(Clk), .Q(Dout[24]), .QN(n32) );
  DF1 Dout_reg_31_ ( .D(n63), .C(Clk), .Q(Dout[31]), .QN(n57) );
  DF3 Dout_reg_28_ ( .D(n66), .C(Clk), .Q(Dout[28]), .QN(n51) );
  DF3 Dout_reg_25_ ( .D(n69), .C(Clk), .Q(Dout[25]), .QN(n35) );
  DF3 Dout_reg_17_ ( .D(n77), .C(Clk), .Q(Dout[17]), .QN(n18) );
  DF1 Dout_reg_26_ ( .D(n68), .C(Clk), .Q(Dout[26]), .QN(n47) );
  INV4 U35 ( .A(Din[28]), .Q(n370) );
  CLKIN4 U36 ( .A(Din[31]), .Q(n367) );
  INV4 U37 ( .A(Din[26]), .Q(n372) );
  INV4 U38 ( .A(Din[30]), .Q(n368) );
  INV3 U39 ( .A(Din[21]), .Q(n375) );
  INV3 U40 ( .A(Din[18]), .Q(n380) );
  INV3 U41 ( .A(Din[27]), .Q(n371) );
  INV3 U42 ( .A(Din[22]), .Q(n377) );
  INV4 U43 ( .A(Din[29]), .Q(n369) );
  CLKIN3 U44 ( .A(Din[16]), .Q(n382) );
  INV3 U45 ( .A(Din[13]), .Q(n385) );
  INV3 U46 ( .A(Din[14]), .Q(n383) );
  CLKIN3 U47 ( .A(Din[8]), .Q(n392) );
  INV3 U48 ( .A(Din[15]), .Q(n384) );
  CLKIN3 U49 ( .A(Din[6]), .Q(n390) );
  INV2 U50 ( .A(Din[25]), .Q(n373) );
  INV2 U51 ( .A(Din[23]), .Q(n376) );
  INV2 U52 ( .A(Din[20]), .Q(n378) );
  INV2 U53 ( .A(Din[19]), .Q(n379) );
  INV2 U54 ( .A(Din[17]), .Q(n381) );
  INV2 U55 ( .A(Din[24]), .Q(n374) );
  INV2 U56 ( .A(Din[11]), .Q(n387) );
  INV2 U57 ( .A(Din[10]), .Q(n391) );
  INV2 U58 ( .A(Din[7]), .Q(n389) );
  INV2 U59 ( .A(Din[12]), .Q(n386) );
  INV2 U60 ( .A(Din[9]), .Q(n393) );
  NAND22 U61 ( .A(n366), .B(n363), .Q(n364) );
  NAND22 U62 ( .A(n366), .B(n363), .Q(n365) );
  NAND22 U63 ( .A(n366), .B(n363), .Q(n104) );
  INV3 U64 ( .A(Reset), .Q(n366) );
  INV3 U65 ( .A(n105), .Q(n363) );
  INV3 U66 ( .A(Din[4]), .Q(n398) );
  INV3 U67 ( .A(Din[5]), .Q(n388) );
  INV3 U68 ( .A(Din[3]), .Q(n396) );
  INV3 U69 ( .A(Din[1]), .Q(n394) );
  INV3 U70 ( .A(Din[2]), .Q(n397) );
  INV3 U71 ( .A(Din[0]), .Q(n395) );
  NOR21 U72 ( .A(Load), .B(Reset), .Q(n105) );
endmodule


module adder_16_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n421, n422,
         n424, n426, n568, n571, n572, n573, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850;

  OAI212 U77 ( .A(n91), .B(n782), .C(n92), .Q(n90) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U141 ( .A(n140), .B(n782), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n782), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n784), .B(n782), .C(n788), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U189 ( .A(n176), .B(n782), .C(n177), .Q(n175) );
  OAI212 U197 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U395 ( .A(n226), .B(n808), .C(n227), .Q(n225) );
  OAI212 U412 ( .A(n573), .B(n248), .C(n249), .Q(n424) );
  OAI212 U438 ( .A(n129), .B(n782), .C(n130), .Q(n128) );
  OAI212 U452 ( .A(n120), .B(n782), .C(n121), .Q(n119) );
  OAI212 U378 ( .A(n73), .B(n782), .C(n74), .Q(n72) );
  OAI212 U429 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U465 ( .A(n42), .B(n782), .C(n43), .Q(n41) );
  OAI212 U401 ( .A(n113), .B(n152), .C(n114), .Q(n426) );
  OAI212 U489 ( .A(n840), .B(n5), .C(n841), .Q(n56) );
  AOI212 U506 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U387 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U388 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI212 U444 ( .A(n194), .B(n798), .C(n195), .Q(n191) );
  OAI212 U453 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U474 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U475 ( .A(n126), .B(n834), .C(n127), .Q(n123) );
  OAI212 U478 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  XNR22 U374 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR22 U454 ( .A(n14), .B(n108), .Q(SUM[24]) );
  OAI212 U426 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U483 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U461 ( .A(n102), .B(n782), .C(n103), .Q(n101) );
  OAI212 U349 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  AOI212 U360 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U447 ( .A(n82), .B(n782), .C(n83), .Q(n81) );
  OAI212 U408 ( .A(n244), .B(n808), .C(n245), .Q(n243) );
  AOI212 U409 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U419 ( .A(n806), .B(n808), .C(n804), .Q(n232) );
  OAI212 U451 ( .A(n268), .B(n248), .C(n249), .Q(n247) );
  OAI212 U440 ( .A(n197), .B(n808), .C(n198), .Q(n196) );
  OAI212 U441 ( .A(n208), .B(n808), .C(n209), .Q(n207) );
  OAI212 U463 ( .A(n151), .B(n782), .C(n152), .Q(n146) );
  OAI212 U497 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U505 ( .A(n88), .B(n825), .C(n89), .Q(n85) );
  NOR21 U350 ( .A(n173), .B(n176), .Q(n171) );
  NOR22 U351 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR23 U352 ( .A(n137), .B(n144), .Q(n135) );
  BUF15 U353 ( .A(n178), .Q(n782) );
  INV0 U354 ( .A(n162), .Q(n830) );
  NOR21 U355 ( .A(n840), .B(n6), .Q(n55) );
  AOI211 U356 ( .A(n277), .B(n269), .C(n270), .Q(n573) );
  NOR22 U357 ( .A(B[1]), .B(A[1]), .Q(n278) );
  XNR22 U358 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XNR22 U359 ( .A(n12), .B(n90), .Q(SUM[26]) );
  XNR22 U361 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XNR22 U362 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U363 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NOR23 U364 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR21 U365 ( .A(B[29]), .B(A[29]), .Q(n61) );
  XNR21 U366 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XNR21 U367 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NOR21 U368 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR21 U369 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR21 U370 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NAND23 U371 ( .A(n568), .B(n272), .Q(n270) );
  NOR22 U372 ( .A(n271), .B(n274), .Q(n269) );
  NAND23 U373 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U375 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR21 U376 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR23 U377 ( .A(B[14]), .B(A[14]), .Q(n194) );
  XNR21 U379 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XOR21 U380 ( .A(n33), .B(n262), .Q(SUM[5]) );
  XOR21 U381 ( .A(n30), .B(n808), .Q(SUM[8]) );
  CLKIN2 U382 ( .A(n244), .Q(n805) );
  INV3 U383 ( .A(n799), .Q(n781) );
  INV3 U384 ( .A(n220), .Q(n799) );
  CLKIN6 U385 ( .A(n157), .Q(n787) );
  NAND22 U386 ( .A(n157), .B(n19), .Q(n421) );
  NAND24 U389 ( .A(n835), .B(n787), .Q(n422) );
  NAND24 U390 ( .A(n571), .B(n572), .Q(SUM[15]) );
  NOR24 U391 ( .A(n181), .B(n219), .Q(n179) );
  NOR23 U392 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR23 U393 ( .A(B[9]), .B(A[9]), .Q(n241) );
  INV3 U394 ( .A(n230), .Q(n802) );
  NAND22 U396 ( .A(n810), .B(n266), .Q(n34) );
  INV3 U397 ( .A(n204), .Q(n798) );
  INV3 U398 ( .A(n151), .Q(n785) );
  NAND23 U399 ( .A(n785), .B(n122), .Q(n120) );
  NAND21 U400 ( .A(n785), .B(n844), .Q(n140) );
  NOR23 U402 ( .A(n223), .B(n230), .Q(n221) );
  NOR22 U403 ( .A(n79), .B(n88), .Q(n77) );
  INV1 U404 ( .A(n6), .Q(n824) );
  INV1 U405 ( .A(n135), .Q(n833) );
  AOI211 U406 ( .A(n789), .B(n122), .C(n123), .Q(n121) );
  NAND21 U407 ( .A(n59), .B(n848), .Q(n46) );
  NAND24 U410 ( .A(n239), .B(n221), .Q(n219) );
  NOR22 U411 ( .A(n252), .B(n255), .Q(n250) );
  AOI212 U413 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  CLKIN2 U414 ( .A(n187), .Q(n794) );
  NAND21 U415 ( .A(n23), .B(n187), .Q(n571) );
  XNR22 U416 ( .A(n31), .B(n254), .Q(SUM[7]) );
  OAI212 U417 ( .A(n219), .B(n808), .C(n781), .Q(n214) );
  INV6 U418 ( .A(n219), .Q(n801) );
  XNR22 U420 ( .A(n13), .B(n101), .Q(SUM[25]) );
  OAI211 U421 ( .A(n188), .B(n808), .C(n189), .Q(n187) );
  NOR24 U422 ( .A(B[3]), .B(A[3]), .Q(n271) );
  XOR22 U423 ( .A(n22), .B(n782), .Q(SUM[16]) );
  NAND24 U424 ( .A(n421), .B(n422), .Q(SUM[19]) );
  NOR24 U425 ( .A(n185), .B(n194), .Q(n183) );
  NOR24 U427 ( .A(B[15]), .B(A[15]), .Q(n185) );
  XNR22 U428 ( .A(n27), .B(n225), .Q(SUM[11]) );
  AOI212 U430 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  NAND22 U431 ( .A(n135), .B(n115), .Q(n113) );
  NOR23 U432 ( .A(n117), .B(n126), .Q(n115) );
  XNR22 U433 ( .A(n24), .B(n196), .Q(SUM[14]) );
  OAI212 U434 ( .A(n786), .B(n782), .C(n790), .Q(n108) );
  INV1 U435 ( .A(n111), .Q(n786) );
  XNR22 U436 ( .A(n18), .B(n146), .Q(SUM[20]) );
  OAI211 U437 ( .A(n53), .B(n782), .C(n54), .Q(n52) );
  NAND21 U439 ( .A(n111), .B(n55), .Q(n53) );
  XNR22 U442 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U443 ( .A(n29), .B(n243), .Q(SUM[9]) );
  XNR22 U445 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U446 ( .A(n20), .B(n164), .Q(SUM[18]) );
  AOI211 U448 ( .A(n813), .B(n810), .C(n811), .Q(n262) );
  XNR22 U449 ( .A(n26), .B(n214), .Q(SUM[12]) );
  INV8 U450 ( .A(n424), .Q(n808) );
  NAND21 U455 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NOR23 U456 ( .A(n205), .B(n212), .Q(n203) );
  NOR22 U457 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NAND22 U458 ( .A(n111), .B(n97), .Q(n91) );
  NOR24 U459 ( .A(n113), .B(n151), .Q(n111) );
  XNR22 U460 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NAND21 U462 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NOR23 U464 ( .A(n99), .B(n106), .Q(n97) );
  AOI212 U466 ( .A(n813), .B(n258), .C(n259), .Q(n257) );
  INV2 U467 ( .A(n268), .Q(n813) );
  OAI211 U468 ( .A(n274), .B(n818), .C(n275), .Q(n273) );
  INV3 U469 ( .A(n277), .Q(n818) );
  OAI211 U470 ( .A(n64), .B(n782), .C(n65), .Q(n63) );
  NAND21 U471 ( .A(n111), .B(n66), .Q(n64) );
  NAND21 U472 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND21 U473 ( .A(n785), .B(n135), .Q(n129) );
  NOR22 U476 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NAND20 U477 ( .A(A[23]), .B(B[23]), .Q(n118) );
  CLKIN0 U479 ( .A(n112), .Q(n790) );
  AOI210 U480 ( .A(n799), .B(n203), .C(n204), .Q(n198) );
  NAND20 U481 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND20 U482 ( .A(n801), .B(n203), .Q(n197) );
  XOR21 U484 ( .A(n32), .B(n257), .Q(SUM[6]) );
  AOI211 U485 ( .A(n426), .B(n66), .C(n67), .Q(n65) );
  INV0 U486 ( .A(n194), .Q(n793) );
  NAND20 U487 ( .A(n827), .B(n80), .Q(n11) );
  NOR21 U488 ( .A(n61), .B(n70), .Q(n59) );
  CLKIN0 U490 ( .A(n136), .Q(n834) );
  NAND20 U491 ( .A(n839), .B(n71), .Q(n10) );
  NAND20 U492 ( .A(n816), .B(n253), .Q(n31) );
  INV0 U493 ( .A(n223), .Q(n800) );
  INV0 U494 ( .A(n278), .Q(n821) );
  NAND21 U495 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND21 U496 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND22 U498 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND22 U499 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND21 U500 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND21 U501 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND22 U502 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND22 U503 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND22 U504 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NAND21 U507 ( .A(B[1]), .B(A[1]), .Q(n279) );
  INV3 U508 ( .A(n152), .Q(n789) );
  AOI210 U509 ( .A(n112), .B(n97), .C(n98), .Q(n92) );
  AOI210 U510 ( .A(n426), .B(n824), .C(n826), .Q(n74) );
  INV0 U511 ( .A(n5), .Q(n826) );
  NOR22 U512 ( .A(n241), .B(n244), .Q(n239) );
  NOR22 U513 ( .A(n155), .B(n162), .Q(n153) );
  INV0 U514 ( .A(n176), .Q(n783) );
  INV0 U515 ( .A(n255), .Q(n807) );
  NAND20 U516 ( .A(n171), .B(n830), .Q(n158) );
  NAND20 U517 ( .A(n845), .B(n107), .Q(n14) );
  INV0 U518 ( .A(n88), .Q(n828) );
  INV0 U519 ( .A(n252), .Q(n816) );
  INV0 U520 ( .A(n99), .Q(n822) );
  INV0 U521 ( .A(n79), .Q(n827) );
  INV0 U522 ( .A(n173), .Q(n838) );
  NAND20 U523 ( .A(n838), .B(n174), .Q(n21) );
  INV0 U524 ( .A(n137), .Q(n832) );
  INV0 U525 ( .A(n117), .Q(n850) );
  XOR20 U526 ( .A(n281), .B(n37), .Q(SUM[1]) );
  AOI210 U527 ( .A(n60), .B(n848), .C(n847), .Q(n47) );
  NAND20 U528 ( .A(n805), .B(n245), .Q(n30) );
  NAND20 U529 ( .A(n812), .B(n275), .Q(n36) );
  INV0 U530 ( .A(n274), .Q(n812) );
  INV0 U531 ( .A(n260), .Q(n809) );
  XNR20 U532 ( .A(n34), .B(n813), .Q(SUM[4]) );
  NAND20 U533 ( .A(n795), .B(n213), .Q(n26) );
  NAND20 U534 ( .A(n815), .B(n272), .Q(n35) );
  INV0 U535 ( .A(n240), .Q(n804) );
  CLKIN0 U536 ( .A(n97), .Q(n823) );
  AOI210 U537 ( .A(n799), .B(n190), .C(n191), .Q(n189) );
  INV0 U538 ( .A(n70), .Q(n839) );
  INV0 U539 ( .A(n213), .Q(n797) );
  INV0 U540 ( .A(n185), .Q(n792) );
  INV0 U541 ( .A(n241), .Q(n829) );
  INV0 U542 ( .A(n205), .Q(n820) );
  NAND20 U543 ( .A(n800), .B(n224), .Q(n27) );
  NAND20 U544 ( .A(n793), .B(n195), .Q(n24) );
  CLKIN0 U545 ( .A(n144), .Q(n844) );
  INV0 U546 ( .A(n265), .Q(n810) );
  INV0 U547 ( .A(n155), .Q(n836) );
  INV0 U548 ( .A(n266), .Q(n811) );
  NAND21 U549 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND21 U550 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NOR22 U551 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NOR22 U552 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NAND20 U553 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND21 U554 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND20 U555 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U556 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND22 U557 ( .A(n111), .B(n824), .Q(n73) );
  NAND20 U558 ( .A(n111), .B(n44), .Q(n42) );
  NAND22 U559 ( .A(n97), .B(n77), .Q(n6) );
  NOR20 U560 ( .A(n46), .B(n6), .Q(n44) );
  NAND22 U561 ( .A(n171), .B(n153), .Q(n151) );
  AOI211 U562 ( .A(n789), .B(n135), .C(n136), .Q(n130) );
  AOI210 U563 ( .A(n426), .B(n55), .C(n56), .Q(n54) );
  INV3 U564 ( .A(n60), .Q(n841) );
  NAND22 U565 ( .A(n791), .B(n794), .Q(n572) );
  INV3 U566 ( .A(n23), .Q(n791) );
  INV3 U567 ( .A(n19), .Q(n835) );
  NAND21 U568 ( .A(n111), .B(n84), .Q(n82) );
  NAND21 U569 ( .A(n111), .B(n845), .Q(n102) );
  NAND22 U570 ( .A(n203), .B(n183), .Q(n181) );
  NAND22 U571 ( .A(n239), .B(n802), .Q(n226) );
  INV3 U572 ( .A(n239), .Q(n806) );
  NAND22 U573 ( .A(n801), .B(n795), .Q(n208) );
  INV0 U574 ( .A(n172), .Q(n788) );
  INV3 U575 ( .A(n203), .Q(n796) );
  INV3 U576 ( .A(n59), .Q(n840) );
  NAND22 U577 ( .A(n828), .B(n89), .Q(n12) );
  AOI211 U578 ( .A(n112), .B(n84), .C(n85), .Q(n83) );
  INV0 U579 ( .A(n98), .Q(n825) );
  NAND21 U580 ( .A(n801), .B(n190), .Q(n188) );
  NOR21 U581 ( .A(n194), .B(n796), .Q(n190) );
  AOI210 U582 ( .A(n172), .B(n830), .C(n831), .Q(n159) );
  INV3 U583 ( .A(n163), .Q(n831) );
  NAND22 U584 ( .A(n279), .B(n821), .Q(n37) );
  NAND22 U585 ( .A(n783), .B(n177), .Q(n22) );
  XOR21 U586 ( .A(n36), .B(n818), .Q(SUM[2]) );
  NAND22 U587 ( .A(n829), .B(n242), .Q(n29) );
  XNR21 U588 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U589 ( .A(n842), .B(n62), .Q(n9) );
  INV3 U590 ( .A(n61), .Q(n842) );
  NAND22 U591 ( .A(n837), .B(n127), .Q(n16) );
  INV3 U592 ( .A(n126), .Q(n837) );
  NAND22 U593 ( .A(n850), .B(n118), .Q(n15) );
  NAND22 U594 ( .A(n848), .B(n51), .Q(n8) );
  NAND22 U595 ( .A(n820), .B(n206), .Q(n25) );
  NAND22 U596 ( .A(n830), .B(n163), .Q(n20) );
  INV3 U597 ( .A(n171), .Q(n784) );
  NAND22 U598 ( .A(n802), .B(n231), .Q(n28) );
  NAND22 U599 ( .A(n807), .B(n256), .Q(n32) );
  INV3 U600 ( .A(n231), .Q(n803) );
  NAND22 U601 ( .A(n844), .B(n145), .Q(n18) );
  NAND22 U602 ( .A(n822), .B(n100), .Q(n13) );
  NAND22 U603 ( .A(n832), .B(n138), .Q(n17) );
  NOR21 U604 ( .A(n126), .B(n833), .Q(n122) );
  NOR21 U605 ( .A(n88), .B(n823), .Q(n84) );
  NAND22 U606 ( .A(n809), .B(n261), .Q(n33) );
  NOR21 U607 ( .A(n70), .B(n6), .Q(n66) );
  NAND22 U608 ( .A(n836), .B(n156), .Q(n19) );
  NOR21 U609 ( .A(n260), .B(n265), .Q(n258) );
  NAND22 U610 ( .A(n792), .B(n186), .Q(n23) );
  AOI211 U611 ( .A(n426), .B(n845), .C(n846), .Q(n103) );
  INV3 U612 ( .A(n107), .Q(n846) );
  AOI210 U613 ( .A(n426), .B(n44), .C(n45), .Q(n43) );
  INV3 U614 ( .A(n51), .Q(n847) );
  AOI211 U615 ( .A(n789), .B(n844), .C(n843), .Q(n141) );
  INV3 U616 ( .A(n145), .Q(n843) );
  AOI211 U617 ( .A(n799), .B(n795), .C(n797), .Q(n209) );
  INV3 U618 ( .A(n106), .Q(n845) );
  INV3 U619 ( .A(n212), .Q(n795) );
  NAND22 U620 ( .A(n814), .B(n815), .Q(n568) );
  INV3 U621 ( .A(n275), .Q(n814) );
  INV3 U622 ( .A(n271), .Q(n815) );
  NAND22 U623 ( .A(n849), .B(n40), .Q(n7) );
  NAND22 U624 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR22 U625 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR22 U626 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR22 U627 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR22 U628 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR22 U629 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR22 U630 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR22 U631 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR22 U632 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR22 U633 ( .A(A[2]), .B(B[2]), .Q(n274) );
  NOR22 U634 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR22 U635 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR21 U636 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NAND22 U637 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND22 U638 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U639 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U640 ( .A(B[3]), .B(A[3]), .Q(n272) );
  NAND21 U641 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NAND22 U642 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND22 U643 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND22 U644 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND22 U645 ( .A(A[11]), .B(B[11]), .Q(n224) );
  INV3 U646 ( .A(n50), .Q(n848) );
  NOR21 U647 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U648 ( .A(n38), .Q(SUM[0]) );
  NAND20 U649 ( .A(n819), .B(n281), .Q(n38) );
  INV3 U650 ( .A(n280), .Q(n819) );
  NOR20 U651 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U652 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U653 ( .A(n39), .Q(n849) );
  NOR21 U654 ( .A(B[31]), .B(A[31]), .Q(n39) );
  AOI210 U655 ( .A(n240), .B(n802), .C(n803), .Q(n227) );
endmodule


module adder_16 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_16_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_15_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n419, n425,
         n427, n430, n434, n436, n440, n443, n510, n514, n589, n597, n601,
         n605, n678, n679, n756, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n904, n905, n906, n907;

  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U298 ( .A(n419), .B(n257), .C(n256), .Q(n254) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n904), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U522 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U559 ( .A(n137), .B(n145), .C(n138), .Q(n136) );
  OAI212 U366 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U474 ( .A(n155), .B(n163), .C(n156), .Q(n154) );
  OAI212 U505 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  NAND23 U349 ( .A(n857), .B(n875), .Q(n434) );
  NOR23 U350 ( .A(n205), .B(n212), .Q(n203) );
  NOR24 U351 ( .A(A[13]), .B(B[13]), .Q(n205) );
  INV6 U352 ( .A(n97), .Q(n856) );
  NAND22 U353 ( .A(B[12]), .B(A[12]), .Q(n213) );
  NOR23 U354 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NAND22 U355 ( .A(n111), .B(n44), .Q(n42) );
  NAND21 U356 ( .A(n111), .B(n859), .Q(n102) );
  NAND21 U357 ( .A(n111), .B(n84), .Q(n82) );
  INV6 U358 ( .A(n53), .Q(n829) );
  NAND24 U359 ( .A(n111), .B(n55), .Q(n53) );
  CLKIN6 U360 ( .A(n107), .Q(n858) );
  OAI211 U361 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  NOR23 U362 ( .A(A[14]), .B(B[14]), .Q(n194) );
  NAND22 U363 ( .A(n875), .B(n863), .Q(n427) );
  NAND23 U364 ( .A(n427), .B(n141), .Q(n139) );
  INV3 U365 ( .A(n838), .Q(n830) );
  NOR23 U367 ( .A(n194), .B(n185), .Q(n183) );
  NOR23 U368 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND21 U369 ( .A(B[15]), .B(A[15]), .Q(n186) );
  NOR22 U370 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U371 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR23 U372 ( .A(n117), .B(n126), .Q(n115) );
  NAND24 U373 ( .A(n135), .B(n115), .Q(n113) );
  NAND23 U374 ( .A(n183), .B(n203), .Q(n181) );
  AOI211 U375 ( .A(n60), .B(n843), .C(n844), .Q(n47) );
  NOR23 U376 ( .A(A[17]), .B(B[17]), .Q(n173) );
  NOR22 U377 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR23 U378 ( .A(A[27]), .B(B[27]), .Q(n79) );
  NOR21 U379 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR22 U380 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND23 U381 ( .A(n440), .B(n65), .Q(n63) );
  NAND22 U382 ( .A(n597), .B(n177), .Q(n175) );
  NAND22 U383 ( .A(B[24]), .B(A[24]), .Q(n107) );
  NAND22 U384 ( .A(n589), .B(n835), .Q(n146) );
  NAND22 U385 ( .A(B[16]), .B(A[16]), .Q(n177) );
  NAND22 U386 ( .A(n605), .B(n877), .Q(n164) );
  XNR21 U387 ( .A(n16), .B(n128), .Q(SUM[22]) );
  INV2 U388 ( .A(n88), .Q(n853) );
  AOI211 U389 ( .A(n860), .B(n135), .C(n136), .Q(n130) );
  OAI211 U390 ( .A(n194), .B(n880), .C(n195), .Q(n191) );
  NAND23 U391 ( .A(n849), .B(n875), .Q(n440) );
  OAI211 U392 ( .A(n226), .B(n895), .C(n227), .Q(n225) );
  CLKIN3 U393 ( .A(n247), .Q(n895) );
  NAND26 U394 ( .A(n510), .B(n100), .Q(n98) );
  NAND26 U395 ( .A(n834), .B(n80), .Q(n78) );
  CLKIN6 U396 ( .A(n89), .Q(n832) );
  NAND20 U397 ( .A(n853), .B(n89), .Q(n12) );
  NAND22 U398 ( .A(B[26]), .B(A[26]), .Q(n89) );
  NOR24 U399 ( .A(B[22]), .B(A[22]), .Q(n126) );
  INV6 U400 ( .A(n99), .Q(n855) );
  INV2 U401 ( .A(n756), .Q(n868) );
  NAND22 U402 ( .A(n848), .B(n71), .Q(n10) );
  OAI210 U403 ( .A(n137), .B(n145), .C(n138), .Q(n756) );
  INV0 U404 ( .A(n137), .Q(n869) );
  NOR24 U405 ( .A(n181), .B(n219), .Q(n179) );
  NAND20 U406 ( .A(n888), .B(n203), .Q(n197) );
  CLKIN3 U407 ( .A(n203), .Q(n882) );
  NAND22 U408 ( .A(n879), .B(n875), .Q(n597) );
  INV15 U409 ( .A(n837), .Q(n875) );
  INV2 U410 ( .A(n220), .Q(n886) );
  OAI212 U411 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  NAND22 U412 ( .A(A[25]), .B(B[25]), .Q(n100) );
  XNR22 U413 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NOR23 U414 ( .A(n847), .B(n6), .Q(n55) );
  INV0 U415 ( .A(n204), .Q(n880) );
  NOR23 U416 ( .A(n230), .B(n223), .Q(n221) );
  CLKIN6 U417 ( .A(n79), .Q(n833) );
  AOI212 U418 ( .A(n840), .B(n852), .C(n850), .Q(n74) );
  NAND24 U419 ( .A(n829), .B(n830), .Q(n831) );
  NAND24 U420 ( .A(n831), .B(n54), .Q(n52) );
  NAND22 U421 ( .A(n832), .B(n833), .Q(n834) );
  CLKIN6 U422 ( .A(n836), .Q(n838) );
  AOI212 U423 ( .A(n840), .B(n859), .C(n858), .Q(n103) );
  NOR24 U424 ( .A(n46), .B(n6), .Q(n44) );
  NAND23 U425 ( .A(n59), .B(n843), .Q(n46) );
  XNR22 U426 ( .A(n12), .B(n90), .Q(SUM[26]) );
  XNR22 U427 ( .A(n17), .B(n139), .Q(SUM[21]) );
  OAI211 U428 ( .A(n895), .B(n197), .C(n198), .Q(n196) );
  NOR24 U429 ( .A(A[19]), .B(B[19]), .Q(n155) );
  AOI212 U430 ( .A(n840), .B(n97), .C(n98), .Q(n92) );
  CLKIN15 U431 ( .A(n839), .Q(n840) );
  CLKIN1 U432 ( .A(n860), .Q(n835) );
  INV2 U433 ( .A(n840), .Q(n861) );
  AOI212 U434 ( .A(n840), .B(n55), .C(n56), .Q(n54) );
  AOI212 U435 ( .A(n840), .B(n66), .C(n67), .Q(n65) );
  NAND24 U436 ( .A(n43), .B(n443), .Q(n41) );
  AOI212 U437 ( .A(n840), .B(n44), .C(n45), .Q(n43) );
  XNR22 U438 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U439 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NOR24 U440 ( .A(B[11]), .B(A[11]), .Q(n223) );
  INV1 U441 ( .A(n162), .Q(n866) );
  OAI212 U442 ( .A(n838), .B(n129), .C(n130), .Q(n128) );
  NAND22 U443 ( .A(n865), .B(n875), .Q(n601) );
  NAND22 U444 ( .A(B[9]), .B(A[9]), .Q(n242) );
  XNR22 U445 ( .A(n15), .B(n119), .Q(SUM[23]) );
  OAI212 U446 ( .A(n120), .B(n838), .C(n121), .Q(n119) );
  NAND21 U447 ( .A(A[13]), .B(B[13]), .Q(n206) );
  AOI211 U448 ( .A(n860), .B(n873), .C(n874), .Q(n141) );
  NOR23 U449 ( .A(n241), .B(n244), .Q(n239) );
  AOI212 U450 ( .A(n115), .B(n136), .C(n116), .Q(n114) );
  AOI212 U451 ( .A(n183), .B(n204), .C(n184), .Q(n182) );
  CLKIN3 U452 ( .A(n212), .Q(n884) );
  XNR22 U453 ( .A(n8), .B(n52), .Q(SUM[30]) );
  INV6 U454 ( .A(n50), .Q(n843) );
  NOR23 U455 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV6 U456 ( .A(n112), .Q(n839) );
  XNR22 U457 ( .A(n11), .B(n81), .Q(SUM[27]) );
  OAI212 U458 ( .A(n82), .B(n838), .C(n83), .Q(n81) );
  XNR22 U459 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR22 U460 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NAND22 U461 ( .A(n171), .B(n875), .Q(n605) );
  OAI212 U462 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  INV1 U463 ( .A(n60), .Q(n845) );
  NAND21 U464 ( .A(B[29]), .B(A[29]), .Q(n62) );
  OAI211 U465 ( .A(n188), .B(n895), .C(n189), .Q(n187) );
  NOR23 U466 ( .A(B[20]), .B(A[20]), .Q(n144) );
  XNR22 U467 ( .A(n21), .B(n175), .Q(SUM[17]) );
  INV3 U468 ( .A(n140), .Q(n863) );
  NAND22 U469 ( .A(n111), .B(n875), .Q(n430) );
  XNR22 U470 ( .A(n20), .B(n164), .Q(SUM[18]) );
  CLKIN1 U471 ( .A(n135), .Q(n870) );
  NOR23 U472 ( .A(n155), .B(n162), .Q(n153) );
  AOI212 U473 ( .A(n84), .B(n840), .C(n85), .Q(n83) );
  OAI212 U475 ( .A(n173), .B(n177), .C(n174), .Q(n172) );
  XNR22 U476 ( .A(n19), .B(n157), .Q(SUM[19]) );
  OAI212 U477 ( .A(n838), .B(n102), .C(n103), .Q(n101) );
  XNR22 U478 ( .A(n7), .B(n41), .Q(SUM[31]) );
  OAI210 U479 ( .A(n895), .B(n208), .C(n209), .Q(n207) );
  OAI210 U480 ( .A(n892), .B(n895), .C(n893), .Q(n232) );
  OAI210 U481 ( .A(n244), .B(n895), .C(n245), .Q(n243) );
  XOR20 U482 ( .A(n30), .B(n895), .Q(SUM[8]) );
  OAI210 U483 ( .A(n177), .B(n173), .C(n174), .Q(n436) );
  NOR23 U484 ( .A(n70), .B(n6), .Q(n66) );
  NOR24 U485 ( .A(n61), .B(n70), .Q(n59) );
  INV0 U486 ( .A(n70), .Q(n848) );
  NOR24 U487 ( .A(B[28]), .B(A[28]), .Q(n70) );
  OAI212 U488 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  INV0 U489 ( .A(n117), .Q(n872) );
  NOR23 U490 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NAND21 U491 ( .A(B[11]), .B(A[11]), .Q(n224) );
  NAND22 U492 ( .A(A[10]), .B(B[10]), .Q(n231) );
  OAI210 U493 ( .A(n245), .B(n241), .C(n242), .Q(n425) );
  NOR24 U494 ( .A(A[29]), .B(B[29]), .Q(n61) );
  OAI210 U495 ( .A(n219), .B(n895), .C(n220), .Q(n214) );
  NOR24 U496 ( .A(A[25]), .B(B[25]), .Q(n99) );
  NAND23 U497 ( .A(n239), .B(n221), .Q(n219) );
  NAND23 U498 ( .A(A[20]), .B(B[20]), .Q(n145) );
  AOI211 U499 ( .A(n860), .B(n122), .C(n123), .Q(n121) );
  NAND22 U500 ( .A(B[23]), .B(A[23]), .Q(n118) );
  NAND28 U501 ( .A(n97), .B(n77), .Q(n6) );
  NOR24 U502 ( .A(n99), .B(n106), .Q(n97) );
  INV2 U503 ( .A(n152), .Q(n860) );
  INV0 U504 ( .A(n155), .Q(n862) );
  NOR24 U506 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND22 U507 ( .A(B[18]), .B(A[18]), .Q(n163) );
  OAI211 U508 ( .A(n88), .B(n854), .C(n89), .Q(n85) );
  INV3 U509 ( .A(n98), .Q(n854) );
  AOI212 U510 ( .A(n98), .B(n679), .C(n78), .Q(n5) );
  AOI212 U511 ( .A(n98), .B(n679), .C(n78), .Q(n678) );
  OAI212 U512 ( .A(n70), .B(n678), .C(n71), .Q(n67) );
  AOI210 U513 ( .A(n886), .B(n203), .C(n204), .Q(n198) );
  NAND22 U514 ( .A(B[17]), .B(A[17]), .Q(n174) );
  OAI212 U515 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  INV0 U516 ( .A(n185), .Q(n876) );
  OAI212 U517 ( .A(n223), .B(n231), .C(n224), .Q(n222) );
  NOR22 U518 ( .A(A[18]), .B(B[18]), .Q(n162) );
  NOR23 U519 ( .A(n79), .B(n88), .Q(n77) );
  NOR22 U520 ( .A(n79), .B(n88), .Q(n679) );
  INV2 U521 ( .A(n106), .Q(n859) );
  NAND21 U523 ( .A(B[19]), .B(A[19]), .Q(n156) );
  INV0 U524 ( .A(n173), .Q(n878) );
  NAND22 U525 ( .A(n111), .B(n97), .Q(n91) );
  NOR24 U526 ( .A(A[21]), .B(B[21]), .Q(n137) );
  NAND21 U527 ( .A(B[27]), .B(A[27]), .Q(n80) );
  OAI212 U528 ( .A(n5), .B(n847), .C(n845), .Q(n56) );
  NAND20 U529 ( .A(n879), .B(n177), .Q(n22) );
  NAND24 U530 ( .A(n171), .B(n153), .Q(n151) );
  NOR22 U531 ( .A(n176), .B(n173), .Q(n171) );
  NAND22 U532 ( .A(n864), .B(n875), .Q(n589) );
  NOR24 U533 ( .A(n144), .B(n137), .Q(n135) );
  INV2 U534 ( .A(n59), .Q(n847) );
  NAND22 U535 ( .A(B[28]), .B(A[28]), .Q(n71) );
  NAND22 U536 ( .A(A[22]), .B(B[22]), .Q(n127) );
  OAI211 U537 ( .A(n126), .B(n868), .C(n127), .Q(n123) );
  INV0 U538 ( .A(n126), .Q(n871) );
  NAND22 U539 ( .A(B[14]), .B(A[14]), .Q(n195) );
  NAND22 U540 ( .A(n138), .B(n869), .Q(n17) );
  NAND22 U541 ( .A(A[21]), .B(B[21]), .Q(n138) );
  AOI212 U542 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  NAND22 U543 ( .A(n843), .B(n51), .Q(n8) );
  NAND21 U544 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND21 U545 ( .A(n859), .B(n107), .Q(n14) );
  NAND22 U546 ( .A(n871), .B(n127), .Q(n16) );
  NAND22 U547 ( .A(n878), .B(n174), .Q(n21) );
  INV6 U548 ( .A(n178), .Q(n836) );
  CLKIN6 U549 ( .A(n836), .Q(n837) );
  NAND22 U550 ( .A(n111), .B(n66), .Q(n64) );
  NAND22 U551 ( .A(n111), .B(n852), .Q(n73) );
  NOR24 U552 ( .A(n113), .B(n151), .Q(n111) );
  OAI211 U553 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  INV1 U554 ( .A(n252), .Q(n896) );
  NOR23 U555 ( .A(n252), .B(n255), .Q(n250) );
  NAND21 U556 ( .A(n864), .B(n122), .Q(n120) );
  INV3 U557 ( .A(n151), .Q(n864) );
  NAND22 U558 ( .A(n842), .B(n875), .Q(n443) );
  INV2 U560 ( .A(n678), .Q(n850) );
  NAND22 U561 ( .A(n851), .B(n875), .Q(n514) );
  NAND22 U562 ( .A(n864), .B(n873), .Q(n140) );
  INV3 U563 ( .A(n144), .Q(n873) );
  NAND21 U564 ( .A(n864), .B(n135), .Q(n129) );
  INV0 U565 ( .A(n239), .Q(n892) );
  AOI212 U566 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  NOR23 U567 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NAND20 U568 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND22 U569 ( .A(n92), .B(n434), .Q(n90) );
  CLKIN0 U570 ( .A(n436), .Q(n877) );
  CLKIN1 U571 ( .A(n425), .Q(n893) );
  INV1 U572 ( .A(n158), .Q(n865) );
  NAND22 U573 ( .A(A[8]), .B(B[8]), .Q(n245) );
  INV2 U574 ( .A(n73), .Q(n851) );
  INV2 U575 ( .A(n91), .Q(n857) );
  NAND20 U576 ( .A(n171), .B(n866), .Q(n158) );
  AOI210 U577 ( .A(n899), .B(n258), .C(n259), .Q(n257) );
  INV0 U578 ( .A(n230), .Q(n889) );
  INV0 U579 ( .A(n176), .Q(n879) );
  NAND20 U580 ( .A(n902), .B(n261), .Q(n33) );
  NOR20 U581 ( .A(B[6]), .B(A[6]), .Q(n419) );
  NOR20 U582 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND21 U583 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U584 ( .A(n39), .Q(n841) );
  NAND20 U585 ( .A(n896), .B(n253), .Q(n31) );
  NAND22 U586 ( .A(n514), .B(n74), .Q(n72) );
  NAND22 U587 ( .A(n430), .B(n861), .Q(n108) );
  INV3 U588 ( .A(n219), .Q(n888) );
  INV3 U589 ( .A(n42), .Q(n842) );
  NAND22 U590 ( .A(n888), .B(n884), .Q(n208) );
  AOI211 U591 ( .A(n886), .B(n884), .C(n885), .Q(n209) );
  INV3 U592 ( .A(n213), .Q(n885) );
  INV3 U593 ( .A(n6), .Q(n852) );
  INV3 U594 ( .A(n64), .Q(n849) );
  INV3 U595 ( .A(n268), .Q(n899) );
  NAND22 U596 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U597 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U598 ( .A(n88), .B(n856), .Q(n84) );
  NOR21 U599 ( .A(n126), .B(n870), .Q(n122) );
  NAND20 U600 ( .A(n239), .B(n889), .Q(n226) );
  AOI211 U601 ( .A(n425), .B(n889), .C(n890), .Q(n227) );
  INV3 U602 ( .A(n231), .Q(n890) );
  NAND22 U603 ( .A(n888), .B(n190), .Q(n188) );
  AOI210 U604 ( .A(n886), .B(n190), .C(n191), .Q(n189) );
  NOR21 U605 ( .A(n194), .B(n882), .Q(n190) );
  NAND22 U606 ( .A(n858), .B(n855), .Q(n510) );
  INV3 U607 ( .A(n51), .Q(n844) );
  NAND22 U608 ( .A(n601), .B(n159), .Q(n157) );
  AOI210 U609 ( .A(n436), .B(n866), .C(n867), .Q(n159) );
  INV3 U610 ( .A(n163), .Q(n867) );
  INV3 U611 ( .A(n145), .Q(n874) );
  INV3 U612 ( .A(n223), .Q(n887) );
  INV3 U613 ( .A(n241), .Q(n894) );
  INV3 U614 ( .A(n244), .Q(n891) );
  INV3 U615 ( .A(n61), .Q(n846) );
  NAND22 U616 ( .A(n898), .B(n272), .Q(n35) );
  INV3 U617 ( .A(n271), .Q(n898) );
  INV3 U618 ( .A(n260), .Q(n902) );
  INV3 U619 ( .A(n265), .Q(n900) );
  INV3 U620 ( .A(n419), .Q(n897) );
  AOI211 U621 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U622 ( .A(n271), .B(n274), .Q(n269) );
  NOR21 U623 ( .A(n260), .B(n265), .Q(n258) );
  INV3 U624 ( .A(n277), .Q(n904) );
  INV3 U625 ( .A(n274), .Q(n907) );
  INV3 U626 ( .A(n278), .Q(n906) );
  INV3 U627 ( .A(n266), .Q(n901) );
  NOR21 U628 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U629 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND22 U630 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND22 U631 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NOR21 U632 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U633 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U634 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U635 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U636 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U637 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND22 U638 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NOR21 U639 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U640 ( .A(A[0]), .B(B[0]), .Q(n281) );
  INV3 U641 ( .A(n280), .Q(n905) );
  NOR21 U642 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U643 ( .A(n846), .B(n62), .Q(n9) );
  NAND22 U644 ( .A(n841), .B(n40), .Q(n7) );
  NAND20 U645 ( .A(n862), .B(n156), .Q(n19) );
  NAND20 U646 ( .A(n873), .B(n145), .Q(n18) );
  NAND20 U647 ( .A(n100), .B(n855), .Q(n13) );
  NAND20 U648 ( .A(n118), .B(n872), .Q(n15) );
  XNR21 U649 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U650 ( .A(n224), .B(n887), .Q(n27) );
  XNR21 U651 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U652 ( .A(n881), .B(n206), .Q(n25) );
  XNR21 U653 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U654 ( .A(n883), .B(n195), .Q(n24) );
  XNR21 U655 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XNR21 U656 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U657 ( .A(n231), .B(n889), .Q(n28) );
  NAND20 U658 ( .A(n866), .B(n163), .Q(n20) );
  NAND20 U659 ( .A(n80), .B(n833), .Q(n11) );
  XNR21 U660 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U661 ( .A(n884), .B(n213), .Q(n26) );
  XNR21 U662 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U663 ( .A(n876), .B(n186), .Q(n23) );
  XNR21 U664 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U665 ( .A(n894), .B(n242), .Q(n29) );
  NAND20 U666 ( .A(n891), .B(n245), .Q(n30) );
  XNR21 U667 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XNR21 U668 ( .A(n34), .B(n899), .Q(SUM[4]) );
  NAND22 U669 ( .A(n900), .B(n266), .Q(n34) );
  XOR21 U670 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND20 U671 ( .A(n897), .B(n256), .Q(n32) );
  XOR21 U672 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U673 ( .A(n899), .B(n900), .C(n901), .Q(n262) );
  INV3 U674 ( .A(n38), .Q(SUM[0]) );
  NAND22 U675 ( .A(n905), .B(n281), .Q(n38) );
  XOR21 U676 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U677 ( .A(n906), .B(n279), .Q(n37) );
  XOR21 U678 ( .A(n36), .B(n904), .Q(SUM[2]) );
  NAND22 U679 ( .A(n907), .B(n275), .Q(n36) );
  INV0 U680 ( .A(n194), .Q(n883) );
  INV0 U681 ( .A(n205), .Q(n881) );
  XOR21 U682 ( .A(n22), .B(n838), .Q(SUM[16]) );
endmodule


module adder_15 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_15_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_14_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n61, n62,
         n67, n68, n69, n70, n71, n74, n75, n76, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n91, n92, n95, n96, n97, n98, n99, n100, n105, n106,
         n107, n108, n109, n112, n113, n114, n115, n116, n121, n122, n123,
         n124, n125, n126, n127, n130, n131, n132, n135, n136, n141, n142,
         n143, n144, n145, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n163, n164, n165, n166, n167,
         n168, n173, n174, n175, n176, n177, n180, n181, n182, n183, n184,
         n189, n190, n191, n192, n193, n194, n195, n198, n199, n200, n203,
         n204, n209, n210, n211, n212, n213, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n228, n229, n230, n231, n236,
         n237, n238, n241, n242, n244, n245, n246, n247, n248, n249, n250,
         n251, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n265, n266, n267, n268, n269, n408, n483, n549, n550, n623,
         n624, n691, n760, n761, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829;

  OAI212 U10 ( .A(n39), .B(n761), .C(n40), .Q(n38) );
  OAI212 U18 ( .A(n57), .B(n47), .C(n48), .Q(n46) );
  OAI212 U36 ( .A(n59), .B(n761), .C(n60), .Q(n58) );
  OAI212 U60 ( .A(n788), .B(n761), .C(n691), .Q(n76) );
  OAI212 U74 ( .A(n88), .B(n761), .C(n89), .Q(n87) );
  OAI212 U94 ( .A(n113), .B(n105), .C(n106), .Q(n100) );
  AOI212 U116 ( .A(n121), .B(n136), .C(n122), .Q(n116) );
  OAI212 U124 ( .A(n126), .B(n761), .C(n127), .Q(n125) );
  OAI212 U134 ( .A(n802), .B(n761), .C(n800), .Q(n132) );
  OAI212 U160 ( .A(n163), .B(n153), .C(n154), .Q(n152) );
  OAI212 U186 ( .A(n181), .B(n173), .C(n174), .Q(n168) );
  OAI212 U226 ( .A(n809), .B(n768), .C(n806), .Q(n200) );
  OAI212 U247 ( .A(n216), .B(n244), .C(n217), .Q(n215) );
  OAI212 U273 ( .A(n242), .B(n236), .C(n237), .Q(n231) );
  OAI212 U296 ( .A(n250), .B(n765), .C(n251), .Q(n249) );
  OAI212 U303 ( .A(n254), .B(n256), .C(n255), .Q(n253) );
  OAI212 U311 ( .A(n263), .B(n259), .C(n260), .Q(n258) );
  OAI212 U317 ( .A(n262), .B(n764), .C(n263), .Q(n261) );
  OAI212 U324 ( .A(n269), .B(n266), .C(n267), .Q(n265) );
  OAI212 U370 ( .A(n212), .B(n768), .C(n213), .Q(n211) );
  OAI212 U442 ( .A(n194), .B(n768), .C(n195), .Q(n193) );
  OAI212 U415 ( .A(n108), .B(n761), .C(n109), .Q(n107) );
  OAI212 U439 ( .A(n156), .B(n768), .C(n157), .Q(n155) );
  OAI212 U465 ( .A(n54), .B(n781), .C(n57), .Q(n53) );
  OAI212 U383 ( .A(n184), .B(n149), .C(n150), .Q(n148) );
  OAI212 U411 ( .A(n115), .B(n761), .C(n116), .Q(n114) );
  OAI212 U419 ( .A(n145), .B(n141), .C(n142), .Q(n136) );
  OAI212 U431 ( .A(n70), .B(n761), .C(n71), .Q(n69) );
  AOI212 U496 ( .A(n245), .B(n253), .C(n246), .Q(n244) );
  OAI212 U368 ( .A(n225), .B(n821), .C(n228), .Q(n224) );
  OAI212 U437 ( .A(n176), .B(n768), .C(n177), .Q(n175) );
  AOI212 U358 ( .A(n215), .B(n147), .C(n148), .Q(n1) );
  AOI212 U382 ( .A(n231), .B(n218), .C(n219), .Q(n217) );
  OAI212 U384 ( .A(n228), .B(n220), .C(n221), .Q(n219) );
  OAI212 U407 ( .A(n144), .B(n761), .C(n145), .Q(n143) );
  AOI212 U621 ( .A(n787), .B(n795), .C(n786), .Q(n691) );
  OAI212 U403 ( .A(n75), .B(n67), .C(n68), .Q(n62) );
  OAI212 U416 ( .A(n95), .B(n85), .C(n86), .Q(n84) );
  OAI212 U429 ( .A(n92), .B(n791), .C(n95), .Q(n91) );
  OAI212 U337 ( .A(n199), .B(n191), .C(n192), .Q(n190) );
  CLKIN3 U338 ( .A(n231), .Q(n821) );
  NAND21 U339 ( .A(B[12]), .B(A[12]), .Q(n210) );
  NOR24 U340 ( .A(B[12]), .B(A[12]), .Q(n209) );
  XNR22 U341 ( .A(n11), .B(n107), .Q(SUM[24]) );
  XNR22 U342 ( .A(n20), .B(n182), .Q(SUM[15]) );
  XNR22 U343 ( .A(n18), .B(n164), .Q(SUM[17]) );
  NAND21 U344 ( .A(B[8]), .B(A[8]), .Q(n237) );
  NOR22 U345 ( .A(n173), .B(n180), .Q(n167) );
  XOR21 U346 ( .A(n26), .B(n229), .Q(SUM[9]) );
  INV3 U347 ( .A(n61), .Q(n780) );
  AOI211 U348 ( .A(n785), .B(n61), .C(n62), .Q(n60) );
  NAND22 U349 ( .A(A[19]), .B(B[19]), .Q(n145) );
  NAND22 U350 ( .A(n3), .B(n782), .Q(n70) );
  NOR22 U351 ( .A(n236), .B(n241), .Q(n230) );
  NOR22 U352 ( .A(B[22]), .B(A[22]), .Q(n123) );
  NOR23 U353 ( .A(B[14]), .B(A[14]), .Q(n191) );
  INV3 U354 ( .A(n199), .Q(n819) );
  XNR21 U355 ( .A(n28), .B(n766), .Q(SUM[7]) );
  AOI211 U356 ( .A(n766), .B(n822), .C(n820), .Q(n238) );
  XOR21 U357 ( .A(n25), .B(n222), .Q(SUM[10]) );
  AOI211 U359 ( .A(n766), .B(n223), .C(n224), .Q(n222) );
  NOR21 U360 ( .A(n160), .B(n816), .Q(n158) );
  INV2 U361 ( .A(n821), .Q(n760) );
  NOR23 U362 ( .A(B[16]), .B(A[16]), .Q(n173) );
  INV3 U363 ( .A(n244), .Q(n766) );
  NAND22 U364 ( .A(A[23]), .B(B[23]), .Q(n113) );
  AOI212 U365 ( .A(n204), .B(n189), .C(n190), .Q(n184) );
  NAND24 U366 ( .A(n483), .B(n210), .Q(n204) );
  OAI212 U367 ( .A(n97), .B(n761), .C(n98), .Q(n96) );
  BUF15 U369 ( .A(n1), .Q(n761) );
  NAND21 U371 ( .A(n797), .B(n99), .Q(n97) );
  AOI211 U372 ( .A(n766), .B(n230), .C(n760), .Q(n229) );
  OAI212 U373 ( .A(n183), .B(n768), .C(n550), .Q(n182) );
  XNR22 U374 ( .A(n9), .B(n87), .Q(SUM[26]) );
  INV8 U375 ( .A(n215), .Q(n768) );
  NOR22 U376 ( .A(B[15]), .B(A[15]), .Q(n180) );
  INV0 U377 ( .A(n220), .Q(n826) );
  NOR23 U378 ( .A(A[10]), .B(B[10]), .Q(n220) );
  NAND20 U379 ( .A(n815), .B(n181), .Q(n20) );
  INV0 U380 ( .A(n181), .Q(n813) );
  OAI211 U381 ( .A(n160), .B(n814), .C(n163), .Q(n159) );
  INV2 U385 ( .A(n168), .Q(n814) );
  NOR24 U386 ( .A(B[8]), .B(A[8]), .Q(n236) );
  INV1 U387 ( .A(n131), .Q(n798) );
  NAND22 U388 ( .A(A[21]), .B(B[21]), .Q(n131) );
  INV6 U389 ( .A(n183), .Q(n810) );
  NOR22 U390 ( .A(n149), .B(n183), .Q(n147) );
  NAND24 U391 ( .A(n203), .B(n189), .Q(n183) );
  INV2 U392 ( .A(n236), .Q(n829) );
  NOR22 U393 ( .A(A[13]), .B(B[13]), .Q(n198) );
  NAND22 U394 ( .A(n810), .B(n815), .Q(n176) );
  XNR22 U395 ( .A(n6), .B(n58), .Q(SUM[29]) );
  NOR22 U396 ( .A(n153), .B(n160), .Q(n151) );
  XNR22 U397 ( .A(n8), .B(n76), .Q(SUM[27]) );
  NAND21 U398 ( .A(A[22]), .B(B[22]), .Q(n124) );
  NAND21 U399 ( .A(A[27]), .B(B[27]), .Q(n75) );
  OAI212 U400 ( .A(n50), .B(n761), .C(n51), .Q(n49) );
  NOR23 U401 ( .A(n191), .B(n198), .Q(n189) );
  XNR22 U402 ( .A(n21), .B(n193), .Q(SUM[14]) );
  XOR22 U404 ( .A(n16), .B(n761), .Q(SUM[19]) );
  NOR22 U405 ( .A(n67), .B(n74), .Q(n61) );
  NOR21 U406 ( .A(B[27]), .B(A[27]), .Q(n74) );
  NAND22 U408 ( .A(n3), .B(n61), .Q(n59) );
  XNR22 U409 ( .A(n10), .B(n96), .Q(SUM[25]) );
  XNR22 U410 ( .A(n15), .B(n143), .Q(SUM[20]) );
  XNR22 U412 ( .A(n13), .B(n125), .Q(SUM[22]) );
  XNR22 U413 ( .A(n12), .B(n114), .Q(SUM[23]) );
  XNR22 U414 ( .A(n22), .B(n200), .Q(SUM[13]) );
  INV1 U417 ( .A(n230), .Q(n823) );
  OAI211 U418 ( .A(n199), .B(n191), .C(n192), .Q(n549) );
  NAND22 U420 ( .A(n818), .B(n199), .Q(n22) );
  NAND22 U421 ( .A(A[13]), .B(B[13]), .Q(n199) );
  XNR22 U422 ( .A(n5), .B(n49), .Q(SUM[30]) );
  INV2 U423 ( .A(n198), .Q(n818) );
  NAND21 U424 ( .A(n796), .B(n124), .Q(n13) );
  OAI211 U425 ( .A(n131), .B(n123), .C(n124), .Q(n122) );
  INV6 U426 ( .A(n550), .Q(n807) );
  AOI212 U427 ( .A(n204), .B(n189), .C(n549), .Q(n550) );
  XNR22 U428 ( .A(n132), .B(n14), .Q(SUM[21]) );
  AOI211 U430 ( .A(n785), .B(n52), .C(n53), .Q(n51) );
  NOR23 U432 ( .A(n141), .B(n144), .Q(n135) );
  NOR22 U433 ( .A(B[20]), .B(A[20]), .Q(n141) );
  NAND21 U434 ( .A(A[14]), .B(B[14]), .Q(n192) );
  CLKIN3 U435 ( .A(n3), .Q(n788) );
  NAND21 U436 ( .A(n3), .B(n776), .Q(n39) );
  NOR23 U438 ( .A(n81), .B(n115), .Q(n3) );
  NOR22 U440 ( .A(n209), .B(n212), .Q(n203) );
  NAND21 U441 ( .A(A[20]), .B(B[20]), .Q(n142) );
  XNR22 U443 ( .A(n7), .B(n69), .Q(SUM[28]) );
  INV2 U444 ( .A(n191), .Q(n817) );
  OAI211 U445 ( .A(n165), .B(n768), .C(n166), .Q(n164) );
  CLKIN2 U446 ( .A(n167), .Q(n816) );
  NAND20 U447 ( .A(n817), .B(n192), .Q(n21) );
  NAND22 U448 ( .A(n810), .B(n158), .Q(n156) );
  NAND21 U449 ( .A(n23), .B(n211), .Q(n623) );
  NAND21 U450 ( .A(A[10]), .B(B[10]), .Q(n221) );
  INV2 U451 ( .A(n23), .Q(n805) );
  INV0 U452 ( .A(n204), .Q(n806) );
  XOR21 U453 ( .A(n24), .B(n768), .Q(SUM[11]) );
  NAND22 U454 ( .A(A[7]), .B(B[7]), .Q(n242) );
  NOR22 U455 ( .A(B[25]), .B(A[25]), .Q(n92) );
  AOI211 U456 ( .A(n100), .B(n83), .C(n84), .Q(n82) );
  INV1 U457 ( .A(n81), .Q(n787) );
  INV0 U458 ( .A(n212), .Q(n812) );
  NAND21 U459 ( .A(A[25]), .B(B[25]), .Q(n95) );
  NAND22 U460 ( .A(n99), .B(n83), .Q(n81) );
  NAND22 U461 ( .A(n135), .B(n121), .Q(n115) );
  AOI211 U462 ( .A(n168), .B(n151), .C(n152), .Q(n150) );
  NAND20 U463 ( .A(n803), .B(n154), .Q(n17) );
  NAND20 U464 ( .A(n792), .B(n106), .Q(n11) );
  NAND21 U466 ( .A(n779), .B(n68), .Q(n7) );
  NAND20 U467 ( .A(n784), .B(n86), .Q(n9) );
  INV0 U468 ( .A(n130), .Q(n799) );
  INV2 U469 ( .A(n250), .Q(n773) );
  NOR21 U470 ( .A(B[29]), .B(A[29]), .Q(n54) );
  NOR20 U471 ( .A(A[31]), .B(B[31]), .Q(n36) );
  INV3 U472 ( .A(n691), .Q(n785) );
  AOI210 U473 ( .A(n807), .B(n167), .C(n168), .Q(n166) );
  NAND20 U474 ( .A(n810), .B(n167), .Q(n165) );
  NAND20 U475 ( .A(n135), .B(n799), .Q(n126) );
  NAND21 U476 ( .A(n797), .B(n794), .Q(n108) );
  NAND20 U477 ( .A(n61), .B(n45), .Q(n43) );
  NOR22 U478 ( .A(n105), .B(n112), .Q(n99) );
  NAND20 U479 ( .A(n827), .B(n228), .Q(n26) );
  INV0 U480 ( .A(n225), .Q(n827) );
  INV1 U481 ( .A(n62), .Q(n781) );
  INV0 U482 ( .A(n144), .Q(n801) );
  NAND20 U483 ( .A(n812), .B(n213), .Q(n24) );
  INV0 U484 ( .A(n105), .Q(n792) );
  INV0 U485 ( .A(n85), .Q(n784) );
  NOR20 U486 ( .A(n250), .B(n247), .Q(n245) );
  OAI211 U487 ( .A(n251), .B(n247), .C(n248), .Q(n246) );
  INV0 U488 ( .A(n67), .Q(n779) );
  NAND20 U489 ( .A(n790), .B(n95), .Q(n10) );
  INV0 U490 ( .A(n160), .Q(n804) );
  INV0 U491 ( .A(n153), .Q(n803) );
  INV0 U492 ( .A(n241), .Q(n822) );
  NAND20 U493 ( .A(n824), .B(n248), .Q(n29) );
  AOI210 U494 ( .A(n204), .B(n818), .C(n819), .Q(n195) );
  NAND20 U495 ( .A(n808), .B(n210), .Q(n23) );
  CLKIN0 U497 ( .A(n112), .Q(n794) );
  NAND21 U498 ( .A(A[15]), .B(B[15]), .Q(n181) );
  NAND21 U499 ( .A(A[17]), .B(B[17]), .Q(n163) );
  NAND20 U500 ( .A(A[18]), .B(B[18]), .Q(n154) );
  NAND20 U501 ( .A(A[26]), .B(B[26]), .Q(n86) );
  NAND20 U502 ( .A(A[24]), .B(B[24]), .Q(n106) );
  NOR20 U503 ( .A(B[30]), .B(A[30]), .Q(n47) );
  NOR20 U504 ( .A(B[5]), .B(A[5]), .Q(n250) );
  NAND20 U505 ( .A(A[29]), .B(B[29]), .Q(n57) );
  NAND20 U506 ( .A(A[30]), .B(B[30]), .Q(n48) );
  NAND20 U507 ( .A(A[28]), .B(B[28]), .Q(n68) );
  INV3 U508 ( .A(n115), .Q(n797) );
  NAND22 U509 ( .A(n797), .B(n789), .Q(n88) );
  CLKIN3 U510 ( .A(n82), .Q(n786) );
  AOI210 U511 ( .A(n795), .B(n99), .C(n100), .Q(n98) );
  NAND22 U512 ( .A(n623), .B(n624), .Q(SUM[12]) );
  NAND22 U513 ( .A(n805), .B(n767), .Q(n624) );
  NAND22 U514 ( .A(n167), .B(n151), .Q(n149) );
  CLKIN3 U515 ( .A(n116), .Q(n795) );
  INV3 U516 ( .A(n211), .Q(n767) );
  NAND20 U517 ( .A(n3), .B(n52), .Q(n50) );
  NAND22 U518 ( .A(n203), .B(n818), .Q(n194) );
  INV0 U519 ( .A(n136), .Q(n800) );
  INV3 U520 ( .A(n408), .Q(n789) );
  NAND22 U521 ( .A(n790), .B(n99), .Q(n408) );
  INV3 U522 ( .A(n203), .Q(n809) );
  INV3 U523 ( .A(n43), .Q(n776) );
  INV3 U524 ( .A(n253), .Q(n765) );
  INV3 U525 ( .A(n265), .Q(n764) );
  NAND22 U526 ( .A(n801), .B(n145), .Q(n16) );
  NAND22 U527 ( .A(n778), .B(n57), .Q(n6) );
  INV3 U528 ( .A(n54), .Q(n778) );
  NAND22 U529 ( .A(n230), .B(n218), .Q(n216) );
  NOR23 U530 ( .A(n220), .B(n225), .Q(n218) );
  NAND22 U531 ( .A(n794), .B(n113), .Q(n12) );
  XOR21 U532 ( .A(n238), .B(n27), .Q(SUM[8]) );
  NAND20 U533 ( .A(n829), .B(n237), .Q(n27) );
  NAND22 U534 ( .A(n826), .B(n221), .Q(n25) );
  INV3 U535 ( .A(n123), .Q(n796) );
  NAND22 U536 ( .A(n775), .B(n48), .Q(n5) );
  INV3 U537 ( .A(n47), .Q(n775) );
  NAND22 U538 ( .A(n822), .B(n242), .Q(n28) );
  XOR21 U539 ( .A(n765), .B(n30), .Q(SUM[5]) );
  NAND22 U540 ( .A(n773), .B(n251), .Q(n30) );
  XNR21 U541 ( .A(n17), .B(n155), .Q(SUM[18]) );
  NAND22 U542 ( .A(n799), .B(n131), .Q(n14) );
  CLKIN0 U543 ( .A(n135), .Q(n802) );
  NAND22 U544 ( .A(n828), .B(n142), .Q(n15) );
  INV3 U545 ( .A(n141), .Q(n828) );
  NAND22 U546 ( .A(n804), .B(n163), .Q(n18) );
  XNR21 U547 ( .A(n19), .B(n175), .Q(SUM[16]) );
  NAND20 U548 ( .A(n174), .B(n825), .Q(n19) );
  INV3 U549 ( .A(n173), .Q(n825) );
  NAND22 U550 ( .A(n782), .B(n75), .Q(n8) );
  NOR21 U551 ( .A(n85), .B(n92), .Q(n83) );
  NOR21 U552 ( .A(n123), .B(n130), .Q(n121) );
  AOI210 U553 ( .A(n136), .B(n799), .C(n798), .Q(n127) );
  AOI211 U554 ( .A(n807), .B(n158), .C(n159), .Q(n157) );
  AOI211 U555 ( .A(n785), .B(n782), .C(n783), .Q(n71) );
  INV3 U556 ( .A(n75), .Q(n783) );
  AOI210 U557 ( .A(n795), .B(n794), .C(n793), .Q(n109) );
  INV3 U558 ( .A(n113), .Q(n793) );
  AOI210 U559 ( .A(n807), .B(n815), .C(n813), .Q(n177) );
  AOI210 U560 ( .A(n795), .B(n789), .C(n91), .Q(n89) );
  INV0 U561 ( .A(n100), .Q(n791) );
  AOI210 U562 ( .A(n785), .B(n776), .C(n777), .Q(n40) );
  INV3 U563 ( .A(n44), .Q(n777) );
  AOI210 U564 ( .A(n62), .B(n45), .C(n46), .Q(n44) );
  NOR20 U565 ( .A(n225), .B(n823), .Q(n223) );
  INV3 U566 ( .A(n74), .Q(n782) );
  INV3 U567 ( .A(n180), .Q(n815) );
  XNR21 U568 ( .A(n29), .B(n249), .Q(SUM[6]) );
  INV2 U569 ( .A(n247), .Q(n824) );
  INV3 U570 ( .A(n209), .Q(n808) );
  NAND22 U571 ( .A(n811), .B(n808), .Q(n483) );
  INV3 U572 ( .A(n213), .Q(n811) );
  INV3 U573 ( .A(n92), .Q(n790) );
  NOR21 U574 ( .A(n54), .B(n780), .Q(n52) );
  INV3 U575 ( .A(n242), .Q(n820) );
  NOR21 U576 ( .A(n47), .B(n54), .Q(n45) );
  XOR21 U577 ( .A(n31), .B(n256), .Q(SUM[4]) );
  NAND22 U578 ( .A(n772), .B(n255), .Q(n31) );
  INV3 U579 ( .A(n254), .Q(n772) );
  XOR21 U580 ( .A(n33), .B(n764), .Q(SUM[2]) );
  NAND22 U581 ( .A(n770), .B(n263), .Q(n33) );
  INV3 U582 ( .A(n262), .Q(n770) );
  XOR21 U583 ( .A(n269), .B(n34), .Q(SUM[1]) );
  NAND22 U584 ( .A(n769), .B(n267), .Q(n34) );
  INV3 U585 ( .A(n266), .Q(n769) );
  XNR21 U586 ( .A(n32), .B(n261), .Q(SUM[3]) );
  NAND22 U587 ( .A(n771), .B(n260), .Q(n32) );
  INV3 U588 ( .A(n259), .Q(n771) );
  AOI211 U589 ( .A(n265), .B(n257), .C(n258), .Q(n256) );
  NOR21 U590 ( .A(n259), .B(n262), .Q(n257) );
  NOR22 U591 ( .A(B[17]), .B(A[17]), .Q(n160) );
  XNR21 U592 ( .A(n4), .B(n38), .Q(SUM[31]) );
  NAND22 U593 ( .A(n774), .B(n37), .Q(n4) );
  NAND22 U594 ( .A(B[31]), .B(A[31]), .Q(n37) );
  NAND22 U595 ( .A(A[9]), .B(B[9]), .Q(n228) );
  NOR21 U596 ( .A(B[28]), .B(A[28]), .Q(n67) );
  NOR22 U597 ( .A(B[24]), .B(A[24]), .Q(n105) );
  NOR22 U598 ( .A(B[18]), .B(A[18]), .Q(n153) );
  NOR22 U599 ( .A(B[26]), .B(A[26]), .Q(n85) );
  NOR21 U600 ( .A(B[19]), .B(A[19]), .Q(n144) );
  NOR22 U601 ( .A(B[11]), .B(A[11]), .Q(n212) );
  NAND22 U602 ( .A(A[6]), .B(B[6]), .Q(n248) );
  NOR21 U603 ( .A(B[23]), .B(A[23]), .Q(n112) );
  NOR21 U604 ( .A(B[21]), .B(A[21]), .Q(n130) );
  NAND22 U605 ( .A(A[11]), .B(B[11]), .Q(n213) );
  INV3 U606 ( .A(n36), .Q(n774) );
  NAND20 U607 ( .A(A[5]), .B(B[5]), .Q(n251) );
  INV3 U608 ( .A(n35), .Q(SUM[0]) );
  NAND22 U609 ( .A(n763), .B(n269), .Q(n35) );
  INV3 U610 ( .A(n268), .Q(n763) );
  NOR20 U611 ( .A(B[0]), .B(A[0]), .Q(n268) );
  NOR20 U612 ( .A(B[3]), .B(A[3]), .Q(n259) );
  NOR20 U613 ( .A(B[2]), .B(A[2]), .Q(n262) );
  NAND20 U614 ( .A(A[0]), .B(B[0]), .Q(n269) );
  NAND20 U615 ( .A(A[2]), .B(B[2]), .Q(n263) );
  NOR20 U616 ( .A(B[1]), .B(A[1]), .Q(n266) );
  NOR20 U617 ( .A(B[4]), .B(A[4]), .Q(n254) );
  NAND20 U618 ( .A(A[1]), .B(B[1]), .Q(n267) );
  NAND20 U619 ( .A(A[3]), .B(B[3]), .Q(n260) );
  NAND20 U620 ( .A(A[4]), .B(B[4]), .Q(n255) );
  NOR21 U622 ( .A(B[6]), .B(A[6]), .Q(n247) );
  NOR22 U623 ( .A(B[7]), .B(A[7]), .Q(n241) );
  NAND22 U624 ( .A(A[16]), .B(B[16]), .Q(n174) );
  NOR23 U625 ( .A(B[9]), .B(A[9]), .Q(n225) );
endmodule


module adder_14 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_14_DW01_add_2 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_13_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n417, n423,
         n426, n427, n438, n439, n506, n507, n508, n510, n586, n587, n742,
         n743, n746, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n900, n901, n902, n903;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U141 ( .A(n140), .B(n829), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n829), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n893), .B(n829), .C(n891), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U189 ( .A(n176), .B(n829), .C(n177), .Q(n175) );
  OAI212 U197 ( .A(n181), .B(n508), .C(n182), .Q(n180) );
  OAI212 U227 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  OAI212 U233 ( .A(n208), .B(n868), .C(n209), .Q(n207) );
  OAI212 U257 ( .A(n226), .B(n868), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n865), .B(n868), .C(n863), .Q(n232) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n901), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U439 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U430 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U425 ( .A(n241), .B(n245), .C(n242), .Q(n240) );
  AOI212 U519 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U416 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U446 ( .A(n73), .B(n829), .C(n74), .Q(n72) );
  OAI212 U488 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U366 ( .A(n219), .B(n868), .C(n220), .Q(n214) );
  OAI212 U401 ( .A(n244), .B(n868), .C(n245), .Q(n243) );
  OAI212 U409 ( .A(n197), .B(n868), .C(n198), .Q(n196) );
  AOI212 U452 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U667 ( .A(n151), .B(n829), .C(n152), .Q(n146) );
  OAI212 U379 ( .A(n185), .B(n195), .C(n186), .Q(n184) );
  OAI212 U417 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  NOR22 U349 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND22 U350 ( .A(n746), .B(n65), .Q(n63) );
  OAI212 U351 ( .A(n835), .B(n5), .C(n833), .Q(n56) );
  NAND21 U352 ( .A(n862), .B(n203), .Q(n197) );
  NAND22 U353 ( .A(n59), .B(n832), .Q(n46) );
  NOR22 U354 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NAND21 U355 ( .A(n171), .B(n850), .Q(n158) );
  INV2 U356 ( .A(n152), .Q(n853) );
  NAND22 U357 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR24 U358 ( .A(n194), .B(n185), .Q(n183) );
  NOR23 U359 ( .A(A[15]), .B(B[15]), .Q(n185) );
  NOR23 U360 ( .A(A[8]), .B(B[8]), .Q(n244) );
  NOR23 U361 ( .A(n79), .B(n88), .Q(n77) );
  XNR22 U362 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NOR22 U363 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND24 U364 ( .A(B[10]), .B(A[10]), .Q(n231) );
  INV6 U365 ( .A(n220), .Q(n859) );
  NOR24 U367 ( .A(n230), .B(n223), .Q(n221) );
  NOR22 U368 ( .A(n117), .B(n126), .Q(n115) );
  NOR22 U369 ( .A(B[23]), .B(A[23]), .Q(n117) );
  INV3 U370 ( .A(n173), .Q(n892) );
  NOR21 U371 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR21 U372 ( .A(n835), .B(n6), .Q(n55) );
  INV3 U373 ( .A(n137), .Q(n873) );
  XOR21 U374 ( .A(n22), .B(n829), .Q(SUM[16]) );
  NOR21 U375 ( .A(n70), .B(n6), .Q(n66) );
  NOR22 U376 ( .A(A[17]), .B(B[17]), .Q(n173) );
  NOR21 U377 ( .A(n194), .B(n880), .Q(n190) );
  INV3 U378 ( .A(n219), .Q(n862) );
  AOI211 U380 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U381 ( .A(B[29]), .B(A[29]), .Q(n61) );
  INV3 U382 ( .A(n231), .Q(n867) );
  NAND23 U383 ( .A(n828), .B(n92), .Q(n90) );
  NAND22 U384 ( .A(n586), .B(n587), .Q(SUM[17]) );
  XNR21 U385 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR21 U386 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NAND22 U387 ( .A(n506), .B(n507), .Q(SUM[14]) );
  NOR23 U388 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND21 U389 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND21 U390 ( .A(n861), .B(n224), .Q(n27) );
  INV1 U391 ( .A(n204), .Q(n878) );
  BUF12 U392 ( .A(n178), .Q(n829) );
  INV3 U393 ( .A(n829), .Q(n827) );
  NAND21 U394 ( .A(A[15]), .B(B[15]), .Q(n186) );
  INV3 U395 ( .A(n205), .Q(n879) );
  NAND22 U396 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NOR24 U397 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NAND24 U398 ( .A(n203), .B(n183), .Q(n181) );
  NOR23 U399 ( .A(n212), .B(n205), .Q(n203) );
  AOI211 U400 ( .A(n853), .B(n135), .C(n136), .Q(n130) );
  CLKIN4 U402 ( .A(n223), .Q(n861) );
  AOI212 U403 ( .A(n112), .B(n848), .C(n847), .Q(n103) );
  NAND22 U404 ( .A(n111), .B(n848), .Q(n102) );
  OAI211 U405 ( .A(n245), .B(n241), .C(n242), .Q(n417) );
  OAI210 U406 ( .A(n42), .B(n829), .C(n43), .Q(n41) );
  OAI211 U407 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  NAND22 U408 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND21 U410 ( .A(n850), .B(n163), .Q(n20) );
  NAND21 U411 ( .A(B[22]), .B(A[22]), .Q(n127) );
  NAND20 U412 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND23 U413 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND24 U414 ( .A(n825), .B(n83), .Q(n81) );
  NOR24 U415 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NOR23 U418 ( .A(n241), .B(n244), .Q(n239) );
  NAND20 U419 ( .A(n866), .B(n231), .Q(n28) );
  INV1 U420 ( .A(n212), .Q(n896) );
  OAI212 U421 ( .A(n868), .B(n188), .C(n189), .Q(n187) );
  NAND24 U422 ( .A(n438), .B(n439), .Q(SUM[25]) );
  INV3 U423 ( .A(n101), .Q(n846) );
  NOR23 U424 ( .A(B[10]), .B(A[10]), .Q(n230) );
  OAI212 U426 ( .A(n852), .B(n829), .C(n854), .Q(n108) );
  NOR23 U427 ( .A(A[13]), .B(B[13]), .Q(n205) );
  NOR22 U428 ( .A(B[12]), .B(A[12]), .Q(n212) );
  OAI210 U429 ( .A(n88), .B(n843), .C(n89), .Q(n85) );
  NOR21 U431 ( .A(n88), .B(n845), .Q(n84) );
  NAND22 U432 ( .A(n253), .B(n869), .Q(n31) );
  NOR20 U433 ( .A(B[4]), .B(A[4]), .Q(n265) );
  CLKIN4 U434 ( .A(n157), .Q(n849) );
  CLKIN0 U435 ( .A(n176), .Q(n897) );
  CLKIN3 U436 ( .A(n175), .Q(n857) );
  NAND22 U437 ( .A(n823), .B(n824), .Q(n825) );
  INV3 U438 ( .A(n82), .Q(n823) );
  INV2 U440 ( .A(n829), .Q(n824) );
  NAND21 U441 ( .A(n111), .B(n84), .Q(n82) );
  INV2 U442 ( .A(n203), .Q(n880) );
  NAND22 U443 ( .A(n826), .B(n827), .Q(n828) );
  INV3 U444 ( .A(n91), .Q(n826) );
  NAND21 U445 ( .A(n111), .B(n97), .Q(n91) );
  INV1 U447 ( .A(n241), .Q(n870) );
  NOR24 U448 ( .A(n113), .B(n151), .Q(n111) );
  CLKIN3 U449 ( .A(n111), .Q(n852) );
  NAND22 U450 ( .A(n111), .B(n55), .Q(n53) );
  NAND22 U451 ( .A(n111), .B(n66), .Q(n64) );
  NAND22 U453 ( .A(n101), .B(n13), .Q(n438) );
  NAND21 U454 ( .A(n186), .B(n856), .Q(n23) );
  NAND28 U455 ( .A(n239), .B(n221), .Q(n219) );
  XNR22 U456 ( .A(n29), .B(n243), .Q(SUM[9]) );
  INV1 U457 ( .A(n194), .Q(n884) );
  NOR23 U458 ( .A(A[14]), .B(B[14]), .Q(n194) );
  XNR22 U459 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NAND26 U460 ( .A(n171), .B(n153), .Q(n151) );
  NOR23 U461 ( .A(n155), .B(n162), .Q(n153) );
  XNR22 U462 ( .A(n225), .B(n27), .Q(SUM[11]) );
  NAND24 U463 ( .A(n135), .B(n115), .Q(n113) );
  OAI212 U464 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  NOR23 U465 ( .A(B[21]), .B(A[21]), .Q(n137) );
  AOI211 U466 ( .A(n853), .B(n122), .C(n123), .Q(n121) );
  XNR22 U467 ( .A(n23), .B(n187), .Q(SUM[15]) );
  AOI212 U468 ( .A(n240), .B(n221), .C(n222), .Q(n508) );
  NAND24 U469 ( .A(n510), .B(n224), .Q(n222) );
  INV0 U470 ( .A(n99), .Q(n844) );
  NOR23 U471 ( .A(n99), .B(n106), .Q(n97) );
  INV2 U472 ( .A(n5), .Q(n840) );
  OAI210 U473 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  XNR22 U474 ( .A(n18), .B(n146), .Q(SUM[20]) );
  OAI211 U475 ( .A(n53), .B(n829), .C(n54), .Q(n52) );
  XNR22 U476 ( .A(n12), .B(n90), .Q(SUM[26]) );
  AOI211 U477 ( .A(n423), .B(n66), .C(n67), .Q(n65) );
  XNR22 U478 ( .A(n28), .B(n232), .Q(SUM[10]) );
  INV2 U479 ( .A(n230), .Q(n866) );
  OAI211 U480 ( .A(n194), .B(n878), .C(n195), .Q(n191) );
  NAND22 U481 ( .A(A[12]), .B(B[12]), .Q(n213) );
  OAI212 U482 ( .A(n129), .B(n829), .C(n130), .Q(n128) );
  INV2 U483 ( .A(n213), .Q(n894) );
  NAND21 U484 ( .A(n896), .B(n213), .Q(n26) );
  AOI212 U485 ( .A(n183), .B(n204), .C(n184), .Q(n182) );
  NOR24 U486 ( .A(n219), .B(n181), .Q(n179) );
  OAI212 U487 ( .A(n120), .B(n829), .C(n121), .Q(n119) );
  OAI211 U489 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  XNR22 U490 ( .A(n25), .B(n207), .Q(SUM[13]) );
  INV1 U491 ( .A(n88), .Q(n841) );
  NAND22 U492 ( .A(n111), .B(n839), .Q(n73) );
  AOI212 U493 ( .A(n423), .B(n839), .C(n840), .Q(n74) );
  INV2 U494 ( .A(n6), .Q(n839) );
  NAND24 U495 ( .A(n742), .B(n743), .Q(SUM[19]) );
  NAND21 U496 ( .A(B[14]), .B(A[14]), .Q(n195) );
  XNR22 U497 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U498 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR22 U499 ( .A(n20), .B(n164), .Q(SUM[18]) );
  XNR22 U500 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND21 U501 ( .A(B[13]), .B(A[13]), .Q(n206) );
  CLKIN3 U502 ( .A(n97), .Q(n845) );
  OAI211 U503 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NAND20 U504 ( .A(n841), .B(n89), .Q(n12) );
  NOR23 U505 ( .A(n173), .B(n176), .Q(n171) );
  NOR22 U506 ( .A(B[16]), .B(A[16]), .Q(n176) );
  XNR22 U507 ( .A(n16), .B(n128), .Q(SUM[22]) );
  OAI212 U508 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  INV2 U509 ( .A(n59), .Q(n835) );
  NAND24 U510 ( .A(n97), .B(n77), .Q(n6) );
  NOR22 U511 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NAND21 U512 ( .A(n851), .B(n122), .Q(n120) );
  INV2 U513 ( .A(n151), .Q(n851) );
  INV0 U514 ( .A(n117), .Q(n875) );
  INV2 U515 ( .A(n64), .Q(n837) );
  NOR22 U516 ( .A(B[22]), .B(A[22]), .Q(n126) );
  OAI211 U517 ( .A(n102), .B(n829), .C(n103), .Q(n101) );
  CLKIN6 U518 ( .A(n247), .Q(n868) );
  NAND21 U520 ( .A(A[24]), .B(B[24]), .Q(n107) );
  INV2 U521 ( .A(n98), .Q(n843) );
  AOI211 U522 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI211 U523 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NAND21 U524 ( .A(B[11]), .B(A[11]), .Q(n224) );
  INV0 U525 ( .A(n155), .Q(n887) );
  NOR22 U526 ( .A(B[19]), .B(A[19]), .Q(n155) );
  AOI211 U527 ( .A(n859), .B(n203), .C(n204), .Q(n198) );
  AOI211 U528 ( .A(n859), .B(n190), .C(n191), .Q(n189) );
  NAND22 U529 ( .A(n862), .B(n190), .Q(n188) );
  NOR22 U530 ( .A(n137), .B(n144), .Q(n135) );
  NOR21 U531 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND21 U532 ( .A(n885), .B(n127), .Q(n16) );
  OAI210 U533 ( .A(n126), .B(n872), .C(n127), .Q(n123) );
  INV2 U534 ( .A(n26), .Q(n895) );
  NAND22 U535 ( .A(n24), .B(n196), .Q(n506) );
  XOR21 U536 ( .A(n30), .B(n868), .Q(SUM[8]) );
  INV0 U537 ( .A(n244), .Q(n864) );
  NAND20 U538 ( .A(n848), .B(n107), .Q(n14) );
  NAND22 U539 ( .A(n834), .B(n62), .Q(n9) );
  INV0 U540 ( .A(n61), .Q(n834) );
  INV0 U541 ( .A(n162), .Q(n850) );
  NAND20 U542 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND20 U543 ( .A(n851), .B(n135), .Q(n129) );
  INV2 U544 ( .A(n24), .Q(n883) );
  NAND21 U545 ( .A(n26), .B(n214), .Q(n426) );
  NAND22 U546 ( .A(n157), .B(n19), .Q(n742) );
  INV0 U547 ( .A(n172), .Q(n891) );
  NOR20 U548 ( .A(n46), .B(n6), .Q(n44) );
  AOI210 U549 ( .A(n417), .B(n866), .C(n867), .Q(n227) );
  CLKIN0 U550 ( .A(n135), .Q(n874) );
  NAND20 U551 ( .A(n239), .B(n866), .Q(n226) );
  NOR20 U552 ( .A(n252), .B(n255), .Q(n250) );
  NAND20 U553 ( .A(n876), .B(n145), .Q(n18) );
  CLKIN0 U554 ( .A(n417), .Q(n863) );
  CLKIN0 U555 ( .A(n185), .Q(n856) );
  NAND20 U556 ( .A(n844), .B(n100), .Q(n13) );
  NAND20 U557 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NOR21 U558 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND20 U559 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NOR20 U560 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND20 U561 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U562 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U563 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U564 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND20 U565 ( .A(A[4]), .B(B[4]), .Q(n266) );
  INV3 U566 ( .A(n214), .Q(n860) );
  NAND20 U567 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U568 ( .A(n196), .Q(n858) );
  INV3 U569 ( .A(n60), .Q(n833) );
  NAND22 U570 ( .A(n883), .B(n858), .Q(n507) );
  NAND22 U571 ( .A(n842), .B(n846), .Q(n439) );
  INV3 U572 ( .A(n13), .Q(n842) );
  NAND22 U573 ( .A(n849), .B(n886), .Q(n743) );
  INV3 U574 ( .A(n19), .Q(n886) );
  NAND22 U575 ( .A(n175), .B(n21), .Q(n586) );
  NAND22 U576 ( .A(n890), .B(n857), .Q(n587) );
  INV3 U577 ( .A(n21), .Q(n890) );
  NAND22 U578 ( .A(n426), .B(n427), .Q(SUM[12]) );
  NAND22 U579 ( .A(n895), .B(n860), .Q(n427) );
  NAND22 U580 ( .A(n837), .B(n827), .Q(n746) );
  NAND22 U581 ( .A(n862), .B(n896), .Q(n208) );
  NAND22 U582 ( .A(n851), .B(n876), .Q(n140) );
  INV3 U583 ( .A(n239), .Q(n865) );
  AOI211 U584 ( .A(n881), .B(n258), .C(n259), .Q(n257) );
  INV3 U585 ( .A(n268), .Q(n881) );
  INV3 U586 ( .A(n277), .Q(n901) );
  NAND22 U587 ( .A(n864), .B(n245), .Q(n30) );
  XOR21 U588 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U589 ( .A(n881), .B(n888), .C(n889), .Q(n262) );
  NAND22 U590 ( .A(n898), .B(n261), .Q(n33) );
  INV3 U591 ( .A(n266), .Q(n889) );
  INV3 U592 ( .A(n126), .Q(n885) );
  NAND22 U593 ( .A(n836), .B(n71), .Q(n10) );
  INV3 U594 ( .A(n70), .Q(n836) );
  NAND22 U595 ( .A(n832), .B(n51), .Q(n8) );
  XNR21 U596 ( .A(n31), .B(n254), .Q(SUM[7]) );
  INV0 U597 ( .A(n252), .Q(n869) );
  XNR21 U598 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U599 ( .A(n882), .B(n272), .Q(n35) );
  INV3 U600 ( .A(n271), .Q(n882) );
  NAND20 U601 ( .A(n879), .B(n206), .Q(n25) );
  AOI210 U602 ( .A(n172), .B(n850), .C(n855), .Q(n159) );
  INV0 U603 ( .A(n163), .Q(n855) );
  NAND20 U604 ( .A(n897), .B(n177), .Q(n22) );
  AOI210 U605 ( .A(n60), .B(n832), .C(n831), .Q(n47) );
  INV3 U606 ( .A(n51), .Q(n831) );
  NAND22 U607 ( .A(n118), .B(n875), .Q(n15) );
  NAND20 U608 ( .A(n870), .B(n242), .Q(n29) );
  NAND22 U609 ( .A(n838), .B(n80), .Q(n11) );
  INV3 U610 ( .A(n79), .Q(n838) );
  NAND22 U611 ( .A(n258), .B(n250), .Q(n248) );
  NAND20 U612 ( .A(n138), .B(n873), .Q(n17) );
  NOR21 U613 ( .A(n61), .B(n70), .Q(n59) );
  INV0 U614 ( .A(n171), .Q(n893) );
  NOR21 U615 ( .A(n126), .B(n874), .Q(n122) );
  NAND20 U616 ( .A(n892), .B(n174), .Q(n21) );
  AOI211 U617 ( .A(n112), .B(n84), .C(n85), .Q(n83) );
  INV0 U618 ( .A(n136), .Q(n872) );
  NAND20 U619 ( .A(n884), .B(n195), .Q(n24) );
  AOI211 U620 ( .A(n859), .B(n896), .C(n894), .Q(n209) );
  INV3 U621 ( .A(n107), .Q(n847) );
  AOI211 U622 ( .A(n853), .B(n876), .C(n877), .Q(n141) );
  INV3 U623 ( .A(n145), .Q(n877) );
  NAND22 U624 ( .A(n156), .B(n887), .Q(n19) );
  INV3 U625 ( .A(n106), .Q(n848) );
  INV3 U626 ( .A(n144), .Q(n876) );
  NAND22 U627 ( .A(n861), .B(n867), .Q(n510) );
  XOR21 U628 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND22 U629 ( .A(n871), .B(n256), .Q(n32) );
  INV2 U630 ( .A(n255), .Q(n871) );
  INV3 U631 ( .A(n260), .Q(n898) );
  INV3 U632 ( .A(n265), .Q(n888) );
  XNR21 U633 ( .A(n34), .B(n881), .Q(SUM[4]) );
  NAND22 U634 ( .A(n888), .B(n266), .Q(n34) );
  XOR21 U635 ( .A(n36), .B(n901), .Q(SUM[2]) );
  NAND22 U636 ( .A(n903), .B(n275), .Q(n36) );
  INV3 U637 ( .A(n274), .Q(n903) );
  XOR21 U638 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U639 ( .A(n902), .B(n279), .Q(n37) );
  INV3 U640 ( .A(n278), .Q(n902) );
  AOI211 U641 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U642 ( .A(n271), .B(n274), .Q(n269) );
  NOR21 U643 ( .A(n260), .B(n265), .Q(n258) );
  XNR21 U644 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U645 ( .A(n830), .B(n40), .Q(n7) );
  NAND20 U646 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV3 U647 ( .A(n50), .Q(n832) );
  NOR20 U648 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U649 ( .A(n39), .Q(n830) );
  NOR20 U650 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND20 U651 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV3 U652 ( .A(n38), .Q(SUM[0]) );
  NAND22 U653 ( .A(n900), .B(n281), .Q(n38) );
  INV3 U654 ( .A(n280), .Q(n900) );
  NOR20 U655 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NOR20 U656 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND20 U657 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U658 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NOR20 U659 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND20 U660 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U661 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NOR20 U662 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NAND21 U663 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND22 U664 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND22 U665 ( .A(A[17]), .B(B[17]), .Q(n174) );
  INV2 U666 ( .A(n112), .Q(n854) );
  AOI210 U668 ( .A(n112), .B(n44), .C(n45), .Q(n43) );
  AOI211 U669 ( .A(n423), .B(n97), .C(n98), .Q(n92) );
  AOI211 U670 ( .A(n423), .B(n55), .C(n56), .Q(n54) );
  OAI212 U671 ( .A(n113), .B(n152), .C(n114), .Q(n423) );
  NAND22 U672 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NOR21 U673 ( .A(B[6]), .B(A[6]), .Q(n255) );
endmodule


module adder_13 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_13_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_12_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n416, n417, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n561, n562, n563, n564,
         n565, n566, n567, n568;

  OAI212 U11 ( .A(n42), .B(n504), .C(n43), .Q(n41) );
  OAI212 U25 ( .A(n53), .B(n505), .C(n54), .Q(n52) );
  OAI212 U39 ( .A(n64), .B(n504), .C(n65), .Q(n63) );
  OAI212 U51 ( .A(n73), .B(n505), .C(n74), .Q(n72) );
  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U65 ( .A(n82), .B(n504), .C(n83), .Q(n81) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n505), .C(n121), .Q(n119) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  AOI212 U195 ( .A(n179), .B(n247), .C(n180), .Q(n178) );
  OAI212 U201 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U207 ( .A(n188), .B(n550), .C(n189), .Q(n187) );
  OAI212 U227 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U329 ( .A(n274), .B(n561), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U496 ( .A(n99), .B(n107), .C(n100), .Q(n98) );
  OAI212 U503 ( .A(n173), .B(n177), .C(n174), .Q(n172) );
  AOI212 U360 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U432 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U392 ( .A(n176), .B(n505), .C(n177), .Q(n175) );
  OAI212 U394 ( .A(n526), .B(n504), .C(n523), .Q(n108) );
  OAI212 U437 ( .A(n129), .B(n505), .C(n130), .Q(n128) );
  OAI212 U445 ( .A(n538), .B(n505), .C(n536), .Q(n164) );
  OAI212 U446 ( .A(n102), .B(n505), .C(n103), .Q(n101) );
  OAI212 U447 ( .A(n504), .B(n140), .C(n141), .Q(n139) );
  OAI212 U452 ( .A(n158), .B(n504), .C(n159), .Q(n157) );
  OAI212 U532 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U534 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U399 ( .A(n208), .B(n550), .C(n209), .Q(n207) );
  OAI212 U522 ( .A(n5), .B(n46), .C(n47), .Q(n45) );
  OAI212 U639 ( .A(n5), .B(n510), .C(n511), .Q(n56) );
  INV3 U349 ( .A(n97), .Q(n519) );
  BUF8 U350 ( .A(B[16]), .Q(n502) );
  NAND21 U351 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NOR23 U352 ( .A(A[17]), .B(B[17]), .Q(n173) );
  NOR24 U353 ( .A(B[6]), .B(A[6]), .Q(n255) );
  INV6 U354 ( .A(n247), .Q(n550) );
  NAND22 U355 ( .A(B[24]), .B(A[24]), .Q(n107) );
  NAND24 U356 ( .A(n135), .B(n417), .Q(n113) );
  CLKIN2 U357 ( .A(n5), .Q(n513) );
  NOR23 U358 ( .A(n99), .B(n106), .Q(n97) );
  NAND22 U359 ( .A(n203), .B(n183), .Q(n181) );
  NOR23 U361 ( .A(n185), .B(n194), .Q(n183) );
  NOR23 U362 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR24 U363 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND22 U364 ( .A(A[25]), .B(B[25]), .Q(n100) );
  AOI212 U365 ( .A(n501), .B(n66), .C(n67), .Q(n65) );
  NAND26 U366 ( .A(n59), .B(n507), .Q(n46) );
  INV2 U367 ( .A(n152), .Q(n531) );
  NOR24 U368 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR24 U369 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NOR22 U370 ( .A(n173), .B(n176), .Q(n171) );
  NOR24 U371 ( .A(n502), .B(n499), .Q(n176) );
  INV1 U372 ( .A(n144), .Q(n529) );
  NOR23 U373 ( .A(B[20]), .B(A[20]), .Q(n144) );
  INV0 U374 ( .A(n70), .Q(n512) );
  NOR21 U375 ( .A(n70), .B(n6), .Q(n66) );
  NOR24 U376 ( .A(n61), .B(n70), .Q(n59) );
  NAND24 U377 ( .A(n171), .B(n153), .Q(n151) );
  NAND26 U378 ( .A(n97), .B(n77), .Q(n6) );
  INV12 U379 ( .A(n503), .Q(n505) );
  NAND22 U380 ( .A(A[14]), .B(B[14]), .Q(n195) );
  INV12 U381 ( .A(n503), .Q(n504) );
  NOR23 U382 ( .A(n155), .B(n162), .Q(n153) );
  NOR23 U383 ( .A(n79), .B(n88), .Q(n77) );
  NOR23 U384 ( .A(n117), .B(n126), .Q(n417) );
  NOR22 U385 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR23 U386 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR23 U387 ( .A(n137), .B(n144), .Q(n135) );
  NOR23 U388 ( .A(B[23]), .B(A[23]), .Q(n117) );
  INV3 U389 ( .A(n59), .Q(n510) );
  NOR23 U390 ( .A(n113), .B(n151), .Q(n111) );
  NOR21 U391 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR21 U393 ( .A(n260), .B(n265), .Q(n258) );
  NOR22 U395 ( .A(n219), .B(n181), .Q(n179) );
  INV3 U396 ( .A(n106), .Q(n520) );
  NOR22 U397 ( .A(A[30]), .B(B[30]), .Q(n50) );
  AOI211 U398 ( .A(n549), .B(n190), .C(n191), .Q(n189) );
  INV2 U400 ( .A(n145), .Q(n530) );
  INV1 U401 ( .A(n137), .Q(n524) );
  NAND26 U402 ( .A(n499), .B(n502), .Q(n177) );
  NAND24 U403 ( .A(B[18]), .B(A[18]), .Q(n163) );
  CLKIN3 U404 ( .A(n61), .Q(n509) );
  INV2 U405 ( .A(n60), .Q(n511) );
  AOI212 U406 ( .A(n60), .B(n507), .C(n508), .Q(n47) );
  XNR22 U407 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND22 U408 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND21 U409 ( .A(n507), .B(n51), .Q(n8) );
  XNR22 U410 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NOR24 U411 ( .A(B[13]), .B(A[13]), .Q(n205) );
  AOI212 U412 ( .A(n501), .B(n84), .C(n85), .Q(n83) );
  XNR22 U413 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NOR24 U414 ( .A(n223), .B(n230), .Q(n221) );
  NAND21 U415 ( .A(A[11]), .B(B[11]), .Q(n224) );
  AOI211 U416 ( .A(n562), .B(n258), .C(n259), .Q(n257) );
  NOR22 U417 ( .A(n241), .B(n244), .Q(n239) );
  CLKIN2 U418 ( .A(n135), .Q(n525) );
  NAND21 U419 ( .A(n533), .B(n135), .Q(n129) );
  INV1 U420 ( .A(n98), .Q(n517) );
  INV1 U421 ( .A(n136), .Q(n522) );
  NAND22 U422 ( .A(A[8]), .B(B[8]), .Q(n245) );
  OAI212 U423 ( .A(n5), .B(n70), .C(n71), .Q(n67) );
  XNR22 U424 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND21 U425 ( .A(B[9]), .B(A[9]), .Q(n242) );
  NAND22 U426 ( .A(n111), .B(n84), .Q(n82) );
  NOR21 U427 ( .A(n88), .B(n519), .Q(n84) );
  XNR22 U428 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U429 ( .A(n20), .B(n164), .Q(SUM[18]) );
  XNR22 U430 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NOR21 U431 ( .A(n126), .B(n525), .Q(n122) );
  AOI212 U433 ( .A(n501), .B(n520), .C(n521), .Q(n103) );
  OAI211 U434 ( .A(n88), .B(n517), .C(n89), .Q(n85) );
  INV0 U435 ( .A(n117), .Q(n527) );
  XNR22 U436 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NOR24 U438 ( .A(B[26]), .B(A[26]), .Q(n88) );
  CLKIN15 U439 ( .A(n500), .Q(n501) );
  XNR22 U440 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NOR23 U441 ( .A(A[18]), .B(B[18]), .Q(n162) );
  NAND22 U442 ( .A(n533), .B(n529), .Q(n140) );
  NAND21 U443 ( .A(A[15]), .B(B[15]), .Q(n186) );
  AOI212 U444 ( .A(n183), .B(n204), .C(n184), .Q(n182) );
  NOR23 U448 ( .A(n252), .B(n255), .Q(n250) );
  XNR22 U449 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NAND21 U450 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND22 U451 ( .A(A[19]), .B(B[19]), .Q(n156) );
  XNR22 U453 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U454 ( .A(n41), .B(n7), .Q(SUM[31]) );
  XNR22 U455 ( .A(n17), .B(n139), .Q(SUM[21]) );
  AOI211 U456 ( .A(n501), .B(n97), .C(n98), .Q(n92) );
  AOI212 U457 ( .A(n501), .B(n44), .C(n45), .Q(n43) );
  NAND22 U458 ( .A(A[26]), .B(B[26]), .Q(n89) );
  INV6 U459 ( .A(n112), .Q(n500) );
  XNR22 U460 ( .A(n18), .B(n146), .Q(SUM[20]) );
  OAI212 U461 ( .A(n151), .B(n504), .C(n498), .Q(n146) );
  INV1 U462 ( .A(n213), .Q(n545) );
  INV2 U463 ( .A(n204), .Q(n544) );
  NOR23 U464 ( .A(n205), .B(n212), .Q(n203) );
  NOR24 U465 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND22 U466 ( .A(n111), .B(n97), .Q(n91) );
  INV2 U467 ( .A(n549), .Q(n497) );
  INV2 U468 ( .A(n220), .Q(n549) );
  XNR22 U469 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI212 U470 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  INV2 U471 ( .A(n531), .Q(n498) );
  OAI211 U472 ( .A(n126), .B(n522), .C(n127), .Q(n123) );
  NOR24 U473 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NAND21 U474 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND22 U475 ( .A(n111), .B(n66), .Q(n64) );
  NOR23 U476 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND21 U477 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND22 U478 ( .A(B[30]), .B(A[30]), .Q(n51) );
  NAND22 U479 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND24 U480 ( .A(n239), .B(n221), .Q(n219) );
  NAND21 U481 ( .A(n528), .B(n127), .Q(n16) );
  NAND22 U482 ( .A(A[28]), .B(B[28]), .Q(n71) );
  OAI212 U483 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  INV0 U484 ( .A(n126), .Q(n528) );
  NOR20 U485 ( .A(n194), .B(n543), .Q(n190) );
  INV0 U486 ( .A(n194), .Q(n540) );
  OAI210 U487 ( .A(n194), .B(n544), .C(n195), .Q(n191) );
  BUF6 U488 ( .A(A[16]), .Q(n499) );
  NAND22 U489 ( .A(n44), .B(n111), .Q(n42) );
  NOR22 U490 ( .A(n46), .B(n6), .Q(n44) );
  OAI210 U491 ( .A(n219), .B(n550), .C(n497), .Q(n214) );
  OAI211 U492 ( .A(n226), .B(n550), .C(n227), .Q(n225) );
  OAI210 U493 ( .A(n553), .B(n550), .C(n554), .Q(n232) );
  OAI211 U494 ( .A(n197), .B(n550), .C(n198), .Q(n196) );
  XOR20 U495 ( .A(n30), .B(n550), .Q(SUM[8]) );
  INV0 U497 ( .A(n99), .Q(n518) );
  OAI211 U498 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI210 U499 ( .A(n173), .B(n177), .C(n174), .Q(n416) );
  NAND21 U500 ( .A(B[23]), .B(A[23]), .Q(n118) );
  INV0 U501 ( .A(n173), .Q(n537) );
  OAI212 U502 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NAND22 U504 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR24 U505 ( .A(A[21]), .B(B[21]), .Q(n137) );
  AOI210 U506 ( .A(n531), .B(n135), .C(n136), .Q(n130) );
  NAND21 U507 ( .A(A[27]), .B(B[27]), .Q(n80) );
  OAI210 U508 ( .A(n244), .B(n550), .C(n245), .Q(n243) );
  INV0 U509 ( .A(n155), .Q(n532) );
  NOR24 U510 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NAND21 U511 ( .A(A[21]), .B(B[21]), .Q(n138) );
  AOI211 U512 ( .A(n549), .B(n203), .C(n204), .Q(n198) );
  AOI211 U513 ( .A(n549), .B(n546), .C(n545), .Q(n209) );
  AOI212 U514 ( .A(n136), .B(n417), .C(n116), .Q(n114) );
  INV2 U515 ( .A(n162), .Q(n535) );
  OAI212 U516 ( .A(n91), .B(n505), .C(n92), .Q(n90) );
  NAND21 U517 ( .A(n548), .B(n546), .Q(n208) );
  NAND22 U518 ( .A(n548), .B(n190), .Q(n188) );
  INV3 U519 ( .A(n219), .Q(n548) );
  AOI212 U520 ( .A(n501), .B(n55), .C(n56), .Q(n54) );
  NOR22 U521 ( .A(n510), .B(n6), .Q(n55) );
  NAND22 U523 ( .A(n512), .B(n71), .Q(n10) );
  NAND21 U524 ( .A(n520), .B(n107), .Q(n14) );
  NAND22 U525 ( .A(n111), .B(n515), .Q(n73) );
  CLKIN12 U526 ( .A(n178), .Q(n503) );
  INV2 U527 ( .A(n6), .Q(n515) );
  NAND20 U528 ( .A(n548), .B(n203), .Q(n197) );
  NOR22 U529 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND21 U530 ( .A(B[12]), .B(A[12]), .Q(n213) );
  INV2 U531 ( .A(n268), .Q(n562) );
  INV2 U533 ( .A(n51), .Q(n508) );
  INV0 U535 ( .A(n239), .Q(n553) );
  AOI212 U536 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  NAND21 U537 ( .A(n533), .B(n122), .Q(n120) );
  AOI211 U538 ( .A(n531), .B(n122), .C(n123), .Q(n121) );
  AOI211 U539 ( .A(n416), .B(n535), .C(n534), .Q(n159) );
  INV0 U540 ( .A(n212), .Q(n546) );
  INV0 U541 ( .A(n277), .Q(n561) );
  INV0 U542 ( .A(n230), .Q(n556) );
  INV0 U543 ( .A(n244), .Q(n557) );
  INV0 U544 ( .A(n274), .Q(n566) );
  INV0 U545 ( .A(n271), .Q(n565) );
  INV0 U546 ( .A(n255), .Q(n559) );
  INV0 U547 ( .A(n252), .Q(n558) );
  INV0 U548 ( .A(n278), .Q(n564) );
  NAND21 U549 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND21 U550 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NOR22 U551 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NAND21 U552 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U553 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND20 U554 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND21 U555 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U556 ( .A(n39), .Q(n506) );
  NAND21 U557 ( .A(n509), .B(n62), .Q(n9) );
  XOR21 U558 ( .A(n22), .B(n504), .Q(SUM[16]) );
  AOI210 U559 ( .A(n562), .B(n567), .C(n568), .Q(n262) );
  XOR21 U560 ( .A(n32), .B(n257), .Q(SUM[6]) );
  XNR20 U561 ( .A(n34), .B(n562), .Q(SUM[4]) );
  NAND20 U562 ( .A(n564), .B(n279), .Q(n37) );
  NAND22 U563 ( .A(n111), .B(n55), .Q(n53) );
  INV3 U564 ( .A(n151), .Q(n533) );
  INV0 U565 ( .A(n240), .Q(n554) );
  INV3 U566 ( .A(n416), .Q(n536) );
  INV3 U567 ( .A(n203), .Q(n543) );
  NAND22 U568 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U569 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U570 ( .A(n271), .B(n274), .Q(n269) );
  NAND20 U571 ( .A(n239), .B(n556), .Q(n226) );
  AOI210 U572 ( .A(n240), .B(n556), .C(n555), .Q(n227) );
  INV3 U573 ( .A(n231), .Q(n555) );
  INV3 U574 ( .A(n107), .Q(n521) );
  INV3 U575 ( .A(n163), .Q(n534) );
  AOI210 U576 ( .A(n531), .B(n529), .C(n530), .Q(n141) );
  NAND22 U577 ( .A(n551), .B(n261), .Q(n33) );
  INV3 U578 ( .A(n260), .Q(n551) );
  INV3 U579 ( .A(n185), .Q(n541) );
  INV3 U580 ( .A(n265), .Q(n567) );
  INV3 U581 ( .A(n88), .Q(n516) );
  INV3 U582 ( .A(n223), .Q(n547) );
  INV3 U583 ( .A(n205), .Q(n542) );
  INV3 U584 ( .A(n241), .Q(n552) );
  INV3 U585 ( .A(n176), .Q(n539) );
  INV3 U586 ( .A(n266), .Q(n568) );
  NOR21 U587 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U588 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U589 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U590 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR21 U591 ( .A(A[12]), .B(B[12]), .Q(n212) );
  NOR21 U592 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U593 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U594 ( .A(A[4]), .B(B[4]), .Q(n266) );
  INV3 U595 ( .A(n50), .Q(n507) );
  NAND22 U596 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NOR21 U597 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U598 ( .A(n280), .Q(n563) );
  NOR21 U599 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U600 ( .A(n516), .B(n89), .Q(n12) );
  NAND22 U601 ( .A(n506), .B(n40), .Q(n7) );
  NAND20 U602 ( .A(n532), .B(n156), .Q(n19) );
  NAND20 U603 ( .A(n529), .B(n145), .Q(n18) );
  NAND20 U604 ( .A(n174), .B(n537), .Q(n21) );
  NAND20 U605 ( .A(n518), .B(n100), .Q(n13) );
  NAND20 U606 ( .A(n527), .B(n118), .Q(n15) );
  NAND20 U607 ( .A(n539), .B(n177), .Q(n22) );
  XNR21 U608 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U609 ( .A(n540), .B(n195), .Q(n24) );
  XNR21 U610 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U611 ( .A(n542), .B(n206), .Q(n25) );
  XNR21 U612 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U613 ( .A(n547), .B(n224), .Q(n27) );
  XNR21 U614 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U615 ( .A(n556), .B(n231), .Q(n28) );
  NAND20 U616 ( .A(n557), .B(n245), .Q(n30) );
  XNR21 U617 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND22 U618 ( .A(n558), .B(n253), .Q(n31) );
  NAND22 U619 ( .A(n567), .B(n266), .Q(n34) );
  XOR21 U620 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND20 U621 ( .A(n535), .B(n163), .Q(n20) );
  NAND20 U622 ( .A(n514), .B(n80), .Q(n11) );
  NAND20 U623 ( .A(n138), .B(n524), .Q(n17) );
  XNR21 U624 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U625 ( .A(n546), .B(n213), .Q(n26) );
  XNR21 U626 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U627 ( .A(n552), .B(n242), .Q(n29) );
  XNR21 U628 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U629 ( .A(n186), .B(n541), .Q(n23) );
  NAND22 U630 ( .A(n559), .B(n256), .Q(n32) );
  XNR21 U631 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND20 U632 ( .A(n565), .B(n272), .Q(n35) );
  XOR21 U633 ( .A(n281), .B(n37), .Q(SUM[1]) );
  XOR21 U634 ( .A(n36), .B(n561), .Q(SUM[2]) );
  NAND20 U635 ( .A(n566), .B(n275), .Q(n36) );
  INV3 U636 ( .A(n38), .Q(SUM[0]) );
  NAND22 U637 ( .A(n563), .B(n281), .Q(n38) );
  INV1 U638 ( .A(n501), .Q(n523) );
  AOI211 U640 ( .A(n501), .B(n515), .C(n513), .Q(n74) );
  CLKIN0 U641 ( .A(n79), .Q(n514) );
  NAND22 U642 ( .A(n111), .B(n520), .Q(n102) );
  INV2 U643 ( .A(n111), .Q(n526) );
  INV1 U644 ( .A(n171), .Q(n538) );
  NAND21 U645 ( .A(n171), .B(n535), .Q(n158) );
endmodule


module adder_12 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_12_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_11_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n418, n424,
         n425, n428, n429, n432, n433, n509, n510, n513, n514, n517, n518,
         n523, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686;

  OAI212 U11 ( .A(n42), .B(n612), .C(n43), .Q(n41) );
  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U77 ( .A(n91), .B(n611), .C(n92), .Q(n90) );
  OAI212 U101 ( .A(n627), .B(n611), .C(n628), .Q(n108) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U127 ( .A(n129), .B(n611), .C(n130), .Q(n128) );
  OAI212 U141 ( .A(n140), .B(n612), .C(n141), .Q(n139) );
  AOI212 U157 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n611), .C(n159), .Q(n157) );
  OAI212 U197 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U207 ( .A(n188), .B(n678), .C(n189), .Q(n187) );
  OAI212 U219 ( .A(n197), .B(n678), .C(n198), .Q(n196) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U233 ( .A(n208), .B(n678), .C(n209), .Q(n207) );
  OAI212 U257 ( .A(n226), .B(n678), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n638), .B(n678), .C(n640), .Q(n232) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U329 ( .A(n274), .B(n676), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U426 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U441 ( .A(n120), .B(n612), .C(n121), .Q(n119) );
  OAI212 U445 ( .A(n604), .B(n173), .C(n174), .Q(n172) );
  OAI212 U427 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U400 ( .A(n53), .B(n612), .C(n54), .Q(n52) );
  OAI212 U404 ( .A(n82), .B(n612), .C(n83), .Q(n81) );
  OAI212 U381 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U416 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U463 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U392 ( .A(n64), .B(n612), .C(n65), .Q(n63) );
  AOI212 U393 ( .A(n240), .B(n221), .C(n523), .Q(n428) );
  OAI212 U407 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  AOI212 U419 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI212 U462 ( .A(n151), .B(n612), .C(n609), .Q(n146) );
  OAI212 U483 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U389 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI212 U391 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U430 ( .A(n245), .B(n241), .C(n242), .Q(n429) );
  OAI212 U437 ( .A(n219), .B(n678), .C(n428), .Q(n214) );
  OAI212 U438 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  NOR24 U519 ( .A(n678), .B(n635), .Q(n418) );
  NAND20 U349 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NOR21 U350 ( .A(B[27]), .B(A[27]), .Q(n79) );
  INV3 U351 ( .A(n135), .Q(n661) );
  NAND23 U352 ( .A(n203), .B(n183), .Q(n181) );
  NOR23 U353 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR23 U354 ( .A(B[14]), .B(A[14]), .Q(n194) );
  XOR22 U355 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND26 U356 ( .A(n602), .B(n103), .Q(n101) );
  NAND22 U357 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NOR24 U358 ( .A(A[13]), .B(B[13]), .Q(n205) );
  NOR23 U359 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NAND22 U360 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NAND24 U361 ( .A(n424), .B(n425), .Q(SUM[27]) );
  INV6 U362 ( .A(n81), .Q(n618) );
  NAND23 U363 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR22 U364 ( .A(n173), .B(n608), .Q(n171) );
  CLKIN6 U365 ( .A(n607), .Q(n608) );
  NAND24 U366 ( .A(n600), .B(n601), .Q(n602) );
  INV3 U367 ( .A(n102), .Q(n600) );
  CLKIN2 U368 ( .A(n611), .Q(n601) );
  NAND22 U369 ( .A(n111), .B(n625), .Q(n102) );
  NOR22 U370 ( .A(B[18]), .B(A[18]), .Q(n162) );
  INV3 U371 ( .A(n177), .Q(n603) );
  INV6 U372 ( .A(n603), .Q(n604) );
  XNR22 U373 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND21 U374 ( .A(n111), .B(n97), .Q(n91) );
  NAND24 U375 ( .A(n97), .B(n77), .Q(n6) );
  NOR22 U376 ( .A(n99), .B(n106), .Q(n97) );
  NOR23 U377 ( .A(n79), .B(n88), .Q(n77) );
  CLKIN6 U378 ( .A(n112), .Q(n605) );
  INV12 U379 ( .A(n605), .Q(n606) );
  INV3 U380 ( .A(n176), .Q(n607) );
  NOR21 U382 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR21 U383 ( .A(B[28]), .B(A[28]), .Q(n70) );
  XNR21 U384 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NOR22 U385 ( .A(n185), .B(n194), .Q(n183) );
  NOR22 U386 ( .A(n117), .B(n126), .Q(n115) );
  NOR22 U387 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR21 U388 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR22 U390 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR21 U394 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR22 U395 ( .A(n155), .B(n162), .Q(n153) );
  INV3 U396 ( .A(n97), .Q(n622) );
  INV3 U397 ( .A(n98), .Q(n623) );
  INV3 U398 ( .A(n151), .Q(n649) );
  NOR22 U399 ( .A(n205), .B(n212), .Q(n203) );
  NAND24 U401 ( .A(n171), .B(n153), .Q(n151) );
  NAND22 U402 ( .A(n517), .B(n518), .Q(SUM[17]) );
  XNR21 U403 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NAND22 U405 ( .A(n646), .B(n634), .Q(n514) );
  INV3 U406 ( .A(n271), .Q(n681) );
  INV3 U408 ( .A(n274), .Q(n680) );
  XNR21 U409 ( .A(n26), .B(n214), .Q(SUM[12]) );
  OAI211 U410 ( .A(n194), .B(n636), .C(n195), .Q(n191) );
  AOI211 U411 ( .A(n606), .B(n620), .C(n617), .Q(n74) );
  NAND21 U412 ( .A(B[13]), .B(A[13]), .Q(n206) );
  OAI211 U413 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  NAND21 U414 ( .A(A[6]), .B(B[6]), .Q(n256) );
  INV4 U415 ( .A(n164), .Q(n631) );
  INV0 U417 ( .A(n647), .Q(n609) );
  INV2 U418 ( .A(n152), .Q(n647) );
  NAND21 U420 ( .A(n649), .B(n135), .Q(n129) );
  NAND23 U421 ( .A(n135), .B(n115), .Q(n113) );
  NOR23 U422 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NAND22 U423 ( .A(n19), .B(n157), .Q(n513) );
  NOR21 U424 ( .A(n88), .B(n622), .Q(n84) );
  NOR21 U425 ( .A(n615), .B(n6), .Q(n55) );
  AOI211 U428 ( .A(n677), .B(n682), .C(n683), .Q(n262) );
  NAND21 U429 ( .A(n645), .B(n118), .Q(n15) );
  INV12 U431 ( .A(n610), .Q(n612) );
  NOR22 U432 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR21 U433 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U434 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND22 U435 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND20 U436 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND24 U439 ( .A(n513), .B(n514), .Q(SUM[19]) );
  NAND24 U440 ( .A(n656), .B(n631), .Q(n510) );
  NAND22 U442 ( .A(n59), .B(n643), .Q(n46) );
  INV15 U443 ( .A(n610), .Q(n611) );
  NAND22 U444 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND21 U446 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NOR22 U447 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND20 U448 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND24 U449 ( .A(n509), .B(n510), .Q(SUM[18]) );
  NOR22 U450 ( .A(A[12]), .B(B[12]), .Q(n212) );
  NAND21 U451 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND22 U452 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NOR21 U453 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR23 U454 ( .A(n230), .B(n223), .Q(n221) );
  NAND24 U455 ( .A(n432), .B(n433), .Q(SUM[21]) );
  NOR20 U456 ( .A(B[4]), .B(A[4]), .Q(n265) );
  OAI210 U457 ( .A(n244), .B(n678), .C(n245), .Q(n243) );
  XNR22 U458 ( .A(n25), .B(n207), .Q(SUM[13]) );
  AOI211 U459 ( .A(n647), .B(n122), .C(n123), .Q(n121) );
  XNR22 U460 ( .A(n23), .B(n187), .Q(SUM[15]) );
  INV0 U461 ( .A(n173), .Q(n664) );
  NAND21 U464 ( .A(A[19]), .B(B[19]), .Q(n156) );
  XNR22 U465 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XNR22 U466 ( .A(n14), .B(n108), .Q(SUM[24]) );
  INV0 U467 ( .A(n205), .Q(n629) );
  NOR22 U468 ( .A(B[23]), .B(A[23]), .Q(n117) );
  OAI212 U469 ( .A(n223), .B(n231), .C(n224), .Q(n222) );
  INV1 U470 ( .A(n241), .Q(n662) );
  NAND21 U471 ( .A(A[17]), .B(B[17]), .Q(n174) );
  XNR22 U472 ( .A(n12), .B(n90), .Q(SUM[26]) );
  XNR22 U473 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NOR20 U474 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR20 U475 ( .A(n271), .B(n274), .Q(n269) );
  OAI210 U476 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  XNR22 U477 ( .A(n15), .B(n119), .Q(SUM[23]) );
  AOI212 U478 ( .A(n606), .B(n625), .C(n624), .Q(n103) );
  AOI210 U479 ( .A(n606), .B(n55), .C(n56), .Q(n54) );
  INV1 U480 ( .A(n88), .Q(n619) );
  INV1 U481 ( .A(n606), .Q(n628) );
  XNR22 U482 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NOR22 U484 ( .A(B[22]), .B(A[22]), .Q(n126) );
  XNR22 U485 ( .A(n13), .B(n101), .Q(SUM[25]) );
  AOI211 U486 ( .A(n606), .B(n97), .C(n98), .Q(n92) );
  AOI211 U487 ( .A(n606), .B(n66), .C(n67), .Q(n65) );
  AOI211 U488 ( .A(n606), .B(n84), .C(n85), .Q(n83) );
  OAI212 U489 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  NAND21 U490 ( .A(n625), .B(n107), .Q(n14) );
  NAND21 U491 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND20 U492 ( .A(n239), .B(n654), .Q(n226) );
  NAND21 U493 ( .A(n231), .B(n654), .Q(n28) );
  INV1 U494 ( .A(n230), .Q(n654) );
  NAND20 U495 ( .A(n667), .B(n604), .Q(n22) );
  OAI212 U496 ( .A(n608), .B(n611), .C(n604), .Q(n175) );
  INV0 U497 ( .A(n223), .Q(n668) );
  OAI211 U498 ( .A(n223), .B(n231), .C(n224), .Q(n523) );
  NAND20 U499 ( .A(A[5]), .B(B[5]), .Q(n261) );
  OAI211 U500 ( .A(n73), .B(n611), .C(n74), .Q(n72) );
  NAND21 U501 ( .A(n111), .B(n55), .Q(n53) );
  CLKIN2 U502 ( .A(n203), .Q(n630) );
  INV3 U503 ( .A(n162), .Q(n657) );
  INV10 U504 ( .A(n178), .Q(n610) );
  OAI210 U505 ( .A(n126), .B(n659), .C(n127), .Q(n123) );
  INV1 U506 ( .A(n126), .Q(n626) );
  CLKIN2 U507 ( .A(n111), .Q(n627) );
  NOR24 U508 ( .A(n113), .B(n151), .Q(n111) );
  INV1 U509 ( .A(n107), .Q(n624) );
  OAI210 U510 ( .A(n88), .B(n623), .C(n89), .Q(n85) );
  NAND21 U511 ( .A(B[11]), .B(A[11]), .Q(n224) );
  INV1 U512 ( .A(n608), .Q(n667) );
  AOI211 U513 ( .A(n641), .B(n203), .C(n204), .Q(n198) );
  INV0 U514 ( .A(n172), .Q(n666) );
  CLKIN0 U515 ( .A(n171), .Q(n665) );
  NAND22 U516 ( .A(n175), .B(n21), .Q(n517) );
  INV2 U517 ( .A(n21), .Q(n663) );
  INV0 U518 ( .A(n163), .Q(n655) );
  NAND21 U520 ( .A(n614), .B(n62), .Q(n9) );
  NAND22 U521 ( .A(n616), .B(n71), .Q(n10) );
  INV0 U522 ( .A(n70), .Q(n616) );
  INV0 U523 ( .A(n144), .Q(n660) );
  CLKIN0 U524 ( .A(n106), .Q(n625) );
  CLKIN0 U525 ( .A(n136), .Q(n659) );
  NAND22 U526 ( .A(n680), .B(n275), .Q(n36) );
  NAND22 U527 ( .A(n681), .B(n272), .Q(n35) );
  INV2 U528 ( .A(n244), .Q(n637) );
  NOR21 U529 ( .A(B[26]), .B(A[26]), .Q(n88) );
  INV1 U530 ( .A(n6), .Q(n620) );
  NOR20 U531 ( .A(n181), .B(n219), .Q(n179) );
  INV2 U532 ( .A(n5), .Q(n617) );
  NOR24 U533 ( .A(n418), .B(n180), .Q(n178) );
  INV2 U534 ( .A(n19), .Q(n646) );
  INV3 U535 ( .A(n428), .Q(n641) );
  CLKIN3 U536 ( .A(n60), .Q(n613) );
  OAI210 U537 ( .A(n615), .B(n5), .C(n613), .Q(n56) );
  NOR20 U538 ( .A(n46), .B(n6), .Q(n44) );
  CLKIN3 U539 ( .A(n59), .Q(n615) );
  CLKIN0 U540 ( .A(n429), .Q(n640) );
  NAND20 U541 ( .A(n239), .B(n221), .Q(n219) );
  NAND20 U542 ( .A(n639), .B(n203), .Q(n197) );
  NAND20 U543 ( .A(n639), .B(n190), .Q(n188) );
  NAND20 U544 ( .A(n639), .B(n652), .Q(n208) );
  XOR20 U545 ( .A(n22), .B(n611), .Q(SUM[16]) );
  INV0 U546 ( .A(n117), .Q(n645) );
  INV0 U547 ( .A(n185), .Q(n650) );
  NAND20 U548 ( .A(n650), .B(n186), .Q(n23) );
  AOI212 U549 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  NAND20 U550 ( .A(n171), .B(n657), .Q(n158) );
  INV0 U551 ( .A(n213), .Q(n651) );
  INV0 U552 ( .A(n61), .Q(n614) );
  NAND20 U553 ( .A(n619), .B(n89), .Q(n12) );
  INV0 U554 ( .A(n99), .Q(n621) );
  NAND21 U555 ( .A(n621), .B(n100), .Q(n13) );
  NAND20 U556 ( .A(n626), .B(n127), .Q(n16) );
  NAND20 U557 ( .A(n662), .B(n242), .Q(n29) );
  NAND20 U558 ( .A(n664), .B(n174), .Q(n21) );
  NAND20 U559 ( .A(n637), .B(n245), .Q(n30) );
  NAND20 U560 ( .A(n657), .B(n163), .Q(n20) );
  INV2 U561 ( .A(n260), .Q(n684) );
  INV0 U562 ( .A(n194), .Q(n673) );
  NAND20 U563 ( .A(n673), .B(n195), .Q(n24) );
  NAND20 U564 ( .A(n652), .B(n213), .Q(n26) );
  INV0 U565 ( .A(n79), .Q(n672) );
  NOR20 U566 ( .A(n241), .B(n244), .Q(n239) );
  NOR20 U567 ( .A(n252), .B(n255), .Q(n250) );
  NOR20 U568 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND20 U569 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U570 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U571 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U572 ( .A(n219), .Q(n639) );
  INV3 U573 ( .A(n179), .Q(n635) );
  INV3 U574 ( .A(n20), .Q(n656) );
  NAND22 U575 ( .A(n669), .B(n632), .Q(n433) );
  INV3 U576 ( .A(n17), .Q(n669) );
  NAND22 U577 ( .A(n633), .B(n663), .Q(n518) );
  NAND22 U578 ( .A(n671), .B(n618), .Q(n425) );
  NAND22 U579 ( .A(n11), .B(n81), .Q(n424) );
  INV3 U580 ( .A(n11), .Q(n671) );
  INV3 U581 ( .A(n139), .Q(n632) );
  INV3 U582 ( .A(n157), .Q(n634) );
  INV3 U583 ( .A(n175), .Q(n633) );
  NAND22 U584 ( .A(n649), .B(n122), .Q(n120) );
  AOI211 U585 ( .A(n677), .B(n258), .C(n259), .Q(n257) );
  INV3 U586 ( .A(n247), .Q(n678) );
  NAND22 U587 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U588 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  INV3 U589 ( .A(n268), .Q(n677) );
  INV3 U590 ( .A(n277), .Q(n676) );
  XNR21 U591 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NOR22 U592 ( .A(n137), .B(n144), .Q(n135) );
  XOR21 U593 ( .A(n30), .B(n678), .Q(SUM[8]) );
  XOR21 U594 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND22 U595 ( .A(n684), .B(n261), .Q(n33) );
  INV3 U596 ( .A(n266), .Q(n683) );
  XOR21 U597 ( .A(n36), .B(n676), .Q(SUM[2]) );
  NAND22 U598 ( .A(n685), .B(n256), .Q(n32) );
  INV3 U599 ( .A(n255), .Q(n685) );
  AOI210 U600 ( .A(n60), .B(n643), .C(n642), .Q(n47) );
  INV3 U601 ( .A(n51), .Q(n642) );
  NAND22 U602 ( .A(n643), .B(n51), .Q(n8) );
  NAND22 U603 ( .A(n660), .B(n145), .Q(n18) );
  NAND22 U604 ( .A(n668), .B(n224), .Q(n27) );
  NAND20 U605 ( .A(n629), .B(n206), .Q(n25) );
  XNR21 U606 ( .A(n34), .B(n677), .Q(SUM[4]) );
  NAND22 U607 ( .A(n682), .B(n266), .Q(n34) );
  XOR21 U608 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U609 ( .A(n679), .B(n279), .Q(n37) );
  INV3 U610 ( .A(n278), .Q(n679) );
  NOR21 U611 ( .A(n61), .B(n70), .Q(n59) );
  NAND22 U612 ( .A(n649), .B(n660), .Q(n140) );
  AOI211 U613 ( .A(n647), .B(n660), .C(n658), .Q(n141) );
  INV3 U614 ( .A(n145), .Q(n658) );
  XNR21 U615 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NOR21 U616 ( .A(n126), .B(n661), .Q(n122) );
  NOR21 U617 ( .A(n194), .B(n630), .Q(n190) );
  XNR21 U618 ( .A(n28), .B(n232), .Q(SUM[10]) );
  INV3 U619 ( .A(n239), .Q(n638) );
  AOI211 U620 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND20 U621 ( .A(n672), .B(n80), .Q(n11) );
  XNR21 U622 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND22 U623 ( .A(n686), .B(n253), .Q(n31) );
  INV3 U624 ( .A(n252), .Q(n686) );
  AOI211 U625 ( .A(n641), .B(n190), .C(n191), .Q(n189) );
  INV0 U626 ( .A(n204), .Q(n636) );
  INV3 U627 ( .A(n265), .Q(n682) );
  AOI211 U628 ( .A(n429), .B(n654), .C(n653), .Q(n227) );
  INV0 U629 ( .A(n231), .Q(n653) );
  AOI211 U630 ( .A(n641), .B(n652), .C(n651), .Q(n209) );
  NAND21 U631 ( .A(n670), .B(n138), .Q(n17) );
  INV0 U632 ( .A(n137), .Q(n670) );
  NOR21 U633 ( .A(n70), .B(n6), .Q(n66) );
  INV3 U634 ( .A(n212), .Q(n652) );
  NAND21 U635 ( .A(n648), .B(n156), .Q(n19) );
  INV0 U636 ( .A(n155), .Q(n648) );
  XNR21 U637 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NOR20 U638 ( .A(n260), .B(n265), .Q(n258) );
  AOI211 U639 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  XNR21 U640 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U641 ( .A(n644), .B(n40), .Q(n7) );
  NAND20 U642 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND22 U643 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND20 U644 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NOR20 U645 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND20 U646 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND21 U647 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND21 U648 ( .A(A[22]), .B(B[22]), .Q(n127) );
  INV3 U649 ( .A(n38), .Q(SUM[0]) );
  NAND22 U650 ( .A(n675), .B(n281), .Q(n38) );
  INV3 U651 ( .A(n280), .Q(n675) );
  NOR20 U652 ( .A(B[0]), .B(A[0]), .Q(n280) );
  INV3 U653 ( .A(n50), .Q(n643) );
  NOR20 U654 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U655 ( .A(n39), .Q(n644) );
  NOR20 U656 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND20 U657 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND20 U658 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U659 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U660 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U661 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U662 ( .A(B[10]), .B(A[10]), .Q(n231) );
  NAND22 U663 ( .A(n111), .B(n84), .Q(n82) );
  NAND22 U664 ( .A(n66), .B(n111), .Q(n64) );
  NAND22 U665 ( .A(n111), .B(n620), .Q(n73) );
  AOI210 U666 ( .A(n647), .B(n135), .C(n136), .Q(n130) );
  NOR22 U667 ( .A(B[21]), .B(A[21]), .Q(n137) );
  OAI212 U668 ( .A(n665), .B(n612), .C(n666), .Q(n164) );
  NOR21 U669 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR21 U670 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND22 U671 ( .A(n17), .B(n139), .Q(n432) );
  NAND22 U672 ( .A(n20), .B(n164), .Q(n509) );
  AOI210 U673 ( .A(n172), .B(n657), .C(n655), .Q(n159) );
  AOI210 U674 ( .A(n606), .B(n44), .C(n45), .Q(n43) );
endmodule


module adder_11 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_11_DW01_add_2 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_10_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n422, n431,
         n432, n434, n439, n440, n443, n444, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n512), .C(n121), .Q(n119) );
  OAI212 U127 ( .A(n129), .B(n512), .C(n130), .Q(n128) );
  OAI212 U141 ( .A(n140), .B(n512), .C(n141), .Q(n139) );
  OAI212 U151 ( .A(n151), .B(n512), .C(n510), .Q(n146) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n512), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n545), .B(n512), .C(n546), .Q(n164) );
  OAI212 U189 ( .A(n176), .B(n512), .C(n177), .Q(n175) );
  OAI212 U227 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U329 ( .A(n274), .B(n560), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U441 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U446 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U448 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U393 ( .A(n241), .B(n245), .C(n242), .Q(n422) );
  OAI222 U397 ( .A(n223), .B(n231), .C(n563), .D(n552), .Q(n222) );
  OAI212 U419 ( .A(n573), .B(n555), .C(n574), .Q(n232) );
  OAI212 U420 ( .A(n244), .B(n555), .C(n245), .Q(n243) );
  OAI212 U421 ( .A(n226), .B(n555), .C(n227), .Q(n225) );
  OAI212 U422 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  XNR22 U485 ( .A(n29), .B(n243), .Q(SUM[9]) );
  OAI212 U486 ( .A(n208), .B(n555), .C(n209), .Q(n207) );
  OAI212 U502 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U404 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  AOI212 U458 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI212 U514 ( .A(n197), .B(n555), .C(n198), .Q(n196) );
  OAI212 U524 ( .A(n188), .B(n555), .C(n189), .Q(n187) );
  OAI212 U643 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  INV2 U349 ( .A(n163), .Q(n538) );
  NOR24 U350 ( .A(A[17]), .B(B[17]), .Q(n173) );
  INV3 U351 ( .A(B[11]), .Q(n552) );
  NOR24 U352 ( .A(n194), .B(n185), .Q(n183) );
  INV2 U353 ( .A(n194), .Q(n550) );
  NOR22 U354 ( .A(n155), .B(n162), .Q(n153) );
  NOR23 U355 ( .A(A[19]), .B(B[19]), .Q(n155) );
  XOR22 U356 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND22 U357 ( .A(n175), .B(n21), .Q(n431) );
  NOR23 U358 ( .A(n205), .B(n212), .Q(n203) );
  CLKIN0 U359 ( .A(n185), .Q(n562) );
  AOI211 U360 ( .A(n422), .B(n221), .C(n222), .Q(n434) );
  NOR24 U361 ( .A(A[11]), .B(B[11]), .Q(n223) );
  NAND21 U362 ( .A(n541), .B(n135), .Q(n129) );
  CLKIN0 U363 ( .A(n135), .Q(n532) );
  NAND23 U364 ( .A(n135), .B(n115), .Q(n113) );
  NAND20 U365 ( .A(B[15]), .B(A[15]), .Q(n186) );
  NAND24 U366 ( .A(n431), .B(n432), .Q(SUM[17]) );
  NAND24 U367 ( .A(n548), .B(n543), .Q(n432) );
  NOR23 U368 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NAND21 U369 ( .A(n111), .B(n66), .Q(n64) );
  NOR22 U370 ( .A(n79), .B(n88), .Q(n77) );
  XNR22 U371 ( .A(n27), .B(n225), .Q(SUM[11]) );
  XNR22 U372 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NOR22 U373 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR23 U374 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND21 U375 ( .A(A[14]), .B(B[14]), .Q(n195) );
  XNR22 U376 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NOR24 U377 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND23 U378 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND22 U379 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND21 U380 ( .A(n554), .B(n203), .Q(n197) );
  INV1 U381 ( .A(n230), .Q(n568) );
  AOI211 U382 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  INV0 U383 ( .A(n231), .Q(n569) );
  NOR21 U384 ( .A(n61), .B(n70), .Q(n59) );
  NOR22 U385 ( .A(n137), .B(n144), .Q(n135) );
  NAND22 U386 ( .A(n97), .B(n77), .Q(n6) );
  INV3 U387 ( .A(n97), .Q(n527) );
  INV3 U388 ( .A(n219), .Q(n554) );
  NAND24 U389 ( .A(n203), .B(n183), .Q(n181) );
  NOR22 U390 ( .A(n173), .B(n176), .Q(n171) );
  NAND22 U391 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND26 U392 ( .A(n239), .B(n221), .Q(n219) );
  NAND23 U394 ( .A(n443), .B(n444), .Q(SUM[21]) );
  NAND22 U395 ( .A(n528), .B(n534), .Q(n444) );
  NAND23 U396 ( .A(n157), .B(n19), .Q(n439) );
  NOR23 U398 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NOR21 U399 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR22 U400 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR24 U401 ( .A(n230), .B(n223), .Q(n221) );
  INV3 U402 ( .A(n112), .Q(n508) );
  INV6 U403 ( .A(n508), .Q(n509) );
  AOI212 U405 ( .A(n509), .B(n84), .C(n85), .Q(n83) );
  CLKIN6 U406 ( .A(n157), .Q(n537) );
  NAND20 U407 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NOR20 U408 ( .A(B[5]), .B(A[5]), .Q(n260) );
  CLKIN0 U409 ( .A(n241), .Q(n579) );
  NAND21 U410 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NOR23 U411 ( .A(B[9]), .B(A[9]), .Q(n241) );
  AOI212 U412 ( .A(n509), .B(n526), .C(n524), .Q(n103) );
  CLKIN4 U413 ( .A(n175), .Q(n548) );
  NOR22 U414 ( .A(B[15]), .B(A[15]), .Q(n185) );
  AOI211 U415 ( .A(n539), .B(n536), .C(n535), .Q(n141) );
  AOI210 U416 ( .A(n539), .B(n135), .C(n136), .Q(n130) );
  INV2 U417 ( .A(n152), .Q(n539) );
  NOR24 U418 ( .A(A[13]), .B(B[13]), .Q(n205) );
  OAI211 U423 ( .A(n53), .B(n512), .C(n54), .Q(n52) );
  AOI210 U424 ( .A(n509), .B(n55), .C(n56), .Q(n54) );
  NOR21 U425 ( .A(n517), .B(n6), .Q(n55) );
  INV2 U426 ( .A(A[11]), .Q(n563) );
  XNR22 U427 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XNR22 U428 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U429 ( .A(A[23]), .B(B[23]), .Q(n118) );
  AOI212 U430 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  CLKIN4 U431 ( .A(n139), .Q(n534) );
  INV2 U432 ( .A(n203), .Q(n566) );
  OAI212 U433 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  NOR23 U434 ( .A(n181), .B(n219), .Q(n179) );
  NAND26 U435 ( .A(n537), .B(n581), .Q(n440) );
  NAND28 U436 ( .A(n439), .B(n440), .Q(SUM[19]) );
  XNR22 U437 ( .A(n26), .B(n214), .Q(SUM[12]) );
  OAI212 U438 ( .A(n219), .B(n555), .C(n434), .Q(n214) );
  BUF15 U439 ( .A(n178), .Q(n512) );
  XNR22 U440 ( .A(n9), .B(n63), .Q(SUM[29]) );
  OAI212 U442 ( .A(n102), .B(n512), .C(n103), .Q(n101) );
  NAND21 U443 ( .A(n111), .B(n526), .Q(n102) );
  XNR22 U444 ( .A(n23), .B(n187), .Q(SUM[15]) );
  XOR21 U445 ( .A(n30), .B(n555), .Q(SUM[8]) );
  NAND21 U447 ( .A(n17), .B(n139), .Q(n443) );
  NOR21 U449 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U450 ( .A(n88), .B(n527), .Q(n84) );
  NOR22 U451 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR22 U452 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NAND21 U453 ( .A(A[21]), .B(B[21]), .Q(n138) );
  INV0 U454 ( .A(n173), .Q(n544) );
  INV1 U455 ( .A(n212), .Q(n577) );
  AOI212 U456 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  NAND20 U457 ( .A(n186), .B(n562), .Q(n23) );
  OAI212 U459 ( .A(n533), .B(n512), .C(n530), .Q(n108) );
  INV1 U460 ( .A(n111), .Q(n533) );
  NAND21 U461 ( .A(n557), .B(n256), .Q(n32) );
  OAI211 U462 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U463 ( .A(n82), .B(n512), .C(n83), .Q(n81) );
  NAND21 U464 ( .A(n111), .B(n84), .Q(n82) );
  NAND22 U465 ( .A(B[12]), .B(A[12]), .Q(n213) );
  OAI211 U466 ( .A(n194), .B(n564), .C(n195), .Q(n191) );
  INV1 U467 ( .A(n539), .Q(n510) );
  OAI212 U468 ( .A(n91), .B(n512), .C(n92), .Q(n90) );
  NAND22 U469 ( .A(A[16]), .B(B[16]), .Q(n177) );
  AOI211 U470 ( .A(n539), .B(n122), .C(n123), .Q(n121) );
  INV1 U471 ( .A(n552), .Q(n511) );
  XNR22 U472 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U473 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI210 U474 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  INV2 U475 ( .A(n5), .Q(n520) );
  OAI210 U476 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  OAI210 U477 ( .A(n88), .B(n525), .C(n89), .Q(n85) );
  XOR21 U478 ( .A(n22), .B(n512), .Q(SUM[16]) );
  XNR22 U479 ( .A(n119), .B(n15), .Q(SUM[23]) );
  XNR22 U480 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NAND21 U481 ( .A(A[26]), .B(B[26]), .Q(n89) );
  XNR22 U482 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U483 ( .A(n20), .B(n164), .Q(SUM[18]) );
  AOI211 U484 ( .A(n551), .B(n190), .C(n191), .Q(n189) );
  NAND21 U487 ( .A(n568), .B(n231), .Q(n28) );
  NAND22 U488 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND21 U489 ( .A(A[20]), .B(B[20]), .Q(n145) );
  OAI212 U490 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  NAND21 U491 ( .A(n536), .B(n145), .Q(n18) );
  INV2 U492 ( .A(n145), .Q(n535) );
  AOI211 U493 ( .A(n509), .B(n97), .C(n98), .Q(n92) );
  INV1 U494 ( .A(n509), .Q(n530) );
  AOI211 U495 ( .A(n509), .B(n66), .C(n67), .Q(n65) );
  INV0 U496 ( .A(n88), .Q(n523) );
  NOR21 U497 ( .A(n126), .B(n532), .Q(n122) );
  XNR22 U498 ( .A(n18), .B(n146), .Q(SUM[20]) );
  OAI212 U499 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  INV0 U500 ( .A(n107), .Q(n524) );
  NAND22 U501 ( .A(n526), .B(n107), .Q(n14) );
  NAND21 U503 ( .A(A[24]), .B(B[24]), .Q(n107) );
  INV3 U504 ( .A(n98), .Q(n525) );
  OAI211 U505 ( .A(n241), .B(n245), .C(n242), .Q(n240) );
  NAND21 U506 ( .A(B[13]), .B(A[13]), .Q(n206) );
  NAND21 U507 ( .A(n577), .B(n213), .Q(n26) );
  INV2 U508 ( .A(n213), .Q(n576) );
  OAI211 U509 ( .A(n73), .B(n512), .C(n74), .Q(n72) );
  OAI211 U510 ( .A(n126), .B(n529), .C(n127), .Q(n123) );
  NAND21 U511 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NOR22 U512 ( .A(n99), .B(n106), .Q(n97) );
  INV0 U513 ( .A(n99), .Q(n583) );
  NOR22 U515 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NAND22 U516 ( .A(n111), .B(n97), .Q(n91) );
  OAI211 U517 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NOR21 U518 ( .A(B[29]), .B(A[29]), .Q(n61) );
  XNR22 U519 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NOR23 U520 ( .A(n113), .B(n151), .Q(n111) );
  INV1 U521 ( .A(n6), .Q(n522) );
  INV2 U522 ( .A(n151), .Q(n541) );
  NOR22 U523 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR21 U525 ( .A(B[28]), .B(A[28]), .Q(n70) );
  INV0 U526 ( .A(n176), .Q(n549) );
  NAND20 U527 ( .A(n239), .B(n568), .Q(n226) );
  CLKIN0 U528 ( .A(n136), .Q(n529) );
  INV0 U529 ( .A(n126), .Q(n547) );
  NAND20 U530 ( .A(n549), .B(n177), .Q(n22) );
  CLKIN0 U531 ( .A(n204), .Q(n564) );
  OAI210 U532 ( .A(n517), .B(n5), .C(n518), .Q(n56) );
  AOI212 U533 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  INV3 U534 ( .A(n434), .Q(n551) );
  NOR20 U535 ( .A(n46), .B(n6), .Q(n44) );
  NOR22 U536 ( .A(n117), .B(n126), .Q(n115) );
  NAND20 U537 ( .A(n516), .B(n62), .Q(n9) );
  NOR20 U538 ( .A(n252), .B(n255), .Q(n250) );
  NAND20 U539 ( .A(n171), .B(n540), .Q(n158) );
  NOR22 U540 ( .A(n241), .B(n244), .Q(n239) );
  INV0 U541 ( .A(n172), .Q(n546) );
  NAND20 U542 ( .A(n540), .B(n163), .Q(n20) );
  NAND20 U543 ( .A(n544), .B(n174), .Q(n21) );
  CLKIN0 U544 ( .A(n244), .Q(n572) );
  NAND21 U545 ( .A(n575), .B(n275), .Q(n36) );
  INV2 U546 ( .A(n274), .Q(n575) );
  INV0 U547 ( .A(n223), .Q(n553) );
  NAND22 U548 ( .A(n553), .B(n224), .Q(n27) );
  CLKIN0 U549 ( .A(n239), .Q(n573) );
  INV0 U550 ( .A(n137), .Q(n531) );
  INV2 U551 ( .A(n260), .Q(n556) );
  CLKIN0 U552 ( .A(n106), .Q(n526) );
  NOR20 U553 ( .A(n260), .B(n265), .Q(n258) );
  NAND21 U554 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND20 U555 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U556 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U557 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U558 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U559 ( .A(n111), .B(n522), .Q(n73) );
  NAND20 U560 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U561 ( .A(n60), .Q(n518) );
  NAND22 U562 ( .A(n171), .B(n153), .Q(n151) );
  AOI211 U563 ( .A(n509), .B(n522), .C(n520), .Q(n74) );
  INV3 U564 ( .A(n19), .Q(n581) );
  INV3 U565 ( .A(n17), .Q(n528) );
  INV3 U566 ( .A(n21), .Q(n543) );
  NAND22 U567 ( .A(n541), .B(n122), .Q(n120) );
  NAND22 U568 ( .A(n554), .B(n190), .Q(n188) );
  NAND22 U569 ( .A(n554), .B(n577), .Q(n208) );
  INV0 U570 ( .A(n422), .Q(n574) );
  INV3 U571 ( .A(n59), .Q(n517) );
  INV3 U572 ( .A(n171), .Q(n545) );
  AOI211 U573 ( .A(n561), .B(n258), .C(n259), .Q(n257) );
  INV3 U574 ( .A(n268), .Q(n561) );
  INV3 U575 ( .A(n277), .Q(n560) );
  NAND22 U576 ( .A(n572), .B(n245), .Q(n30) );
  INV3 U577 ( .A(n255), .Q(n557) );
  XOR21 U578 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U579 ( .A(n561), .B(n570), .C(n571), .Q(n262) );
  NAND22 U580 ( .A(n556), .B(n261), .Q(n33) );
  INV3 U581 ( .A(n266), .Q(n571) );
  NAND22 U582 ( .A(n519), .B(n71), .Q(n10) );
  INV3 U583 ( .A(n70), .Q(n519) );
  NAND22 U584 ( .A(n541), .B(n536), .Q(n140) );
  NAND22 U585 ( .A(n523), .B(n89), .Q(n12) );
  NAND22 U586 ( .A(n521), .B(n80), .Q(n11) );
  INV0 U587 ( .A(n79), .Q(n521) );
  NAND20 U588 ( .A(n542), .B(n118), .Q(n15) );
  INV3 U589 ( .A(n117), .Q(n542) );
  NAND20 U590 ( .A(n195), .B(n550), .Q(n24) );
  NAND20 U591 ( .A(n565), .B(n206), .Q(n25) );
  INV3 U592 ( .A(n205), .Q(n565) );
  NAND22 U593 ( .A(n547), .B(n127), .Q(n16) );
  XNR21 U594 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U595 ( .A(n567), .B(n253), .Q(n31) );
  INV0 U596 ( .A(n252), .Q(n567) );
  XNR21 U597 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND22 U598 ( .A(n515), .B(n51), .Q(n8) );
  NAND20 U599 ( .A(n111), .B(n55), .Q(n53) );
  XOR21 U600 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U601 ( .A(n578), .B(n279), .Q(n37) );
  INV3 U602 ( .A(n278), .Q(n578) );
  NAND20 U603 ( .A(n579), .B(n242), .Q(n29) );
  INV3 U604 ( .A(n61), .Q(n516) );
  AOI210 U605 ( .A(n60), .B(n515), .C(n514), .Q(n47) );
  INV3 U606 ( .A(n51), .Q(n514) );
  NAND20 U607 ( .A(n583), .B(n100), .Q(n13) );
  NAND22 U608 ( .A(n258), .B(n250), .Q(n248) );
  NOR21 U609 ( .A(n194), .B(n566), .Q(n190) );
  NOR21 U610 ( .A(n70), .B(n6), .Q(n66) );
  NAND21 U611 ( .A(n582), .B(n156), .Q(n19) );
  INV0 U612 ( .A(n155), .Q(n582) );
  AOI210 U613 ( .A(n422), .B(n568), .C(n569), .Q(n227) );
  INV3 U614 ( .A(n265), .Q(n570) );
  AOI211 U615 ( .A(n551), .B(n577), .C(n576), .Q(n209) );
  NAND22 U616 ( .A(n531), .B(n138), .Q(n17) );
  NAND20 U617 ( .A(n59), .B(n515), .Q(n46) );
  INV3 U618 ( .A(n144), .Q(n536) );
  INV3 U619 ( .A(n162), .Q(n540) );
  XNR21 U620 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U621 ( .A(n580), .B(n272), .Q(n35) );
  INV2 U622 ( .A(n271), .Q(n580) );
  XNR21 U623 ( .A(n34), .B(n561), .Q(SUM[4]) );
  NAND22 U624 ( .A(n570), .B(n266), .Q(n34) );
  XOR21 U625 ( .A(n36), .B(n560), .Q(SUM[2]) );
  AOI211 U626 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR20 U627 ( .A(n271), .B(n274), .Q(n269) );
  XNR21 U628 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U629 ( .A(n513), .B(n40), .Q(n7) );
  NAND20 U630 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR20 U631 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NOR22 U632 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR22 U633 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR21 U634 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR22 U635 ( .A(B[12]), .B(A[12]), .Q(n212) );
  INV3 U636 ( .A(n50), .Q(n515) );
  NOR20 U637 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND20 U638 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV3 U639 ( .A(n38), .Q(SUM[0]) );
  NAND22 U640 ( .A(n559), .B(n281), .Q(n38) );
  INV3 U641 ( .A(n280), .Q(n559) );
  NOR20 U642 ( .A(B[0]), .B(A[0]), .Q(n280) );
  INV3 U644 ( .A(n39), .Q(n513) );
  NOR20 U645 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND20 U646 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND20 U647 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U648 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U649 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NOR21 U650 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U651 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NAND21 U652 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND21 U653 ( .A(A[19]), .B(B[19]), .Q(n156) );
  AOI210 U654 ( .A(n172), .B(n540), .C(n538), .Q(n159) );
  INV6 U655 ( .A(n247), .Q(n555) );
  NAND21 U656 ( .A(B[17]), .B(A[17]), .Q(n174) );
  NOR22 U657 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND20 U658 ( .A(A[11]), .B(n511), .Q(n224) );
  AOI210 U659 ( .A(n551), .B(n203), .C(n204), .Q(n198) );
  OAI210 U660 ( .A(n42), .B(n512), .C(n43), .Q(n41) );
  OAI211 U661 ( .A(n64), .B(n512), .C(n65), .Q(n63) );
  AOI210 U662 ( .A(n509), .B(n44), .C(n45), .Q(n43) );
endmodule


module adder_10 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_10_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module reg_3 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32,
         n35, n47, n49, n51, n53, n55, n57, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n58, n59, n60, n61, n62, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n104, n105, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395;

  DF3 Dout_reg_16_ ( .D(n78), .C(Clk), .Q(Dout[16]), .QN(n16) );
  DF3 Dout_reg_15_ ( .D(n79), .C(Clk), .Q(Dout[15]), .QN(n14) );
  DF3 Dout_reg_14_ ( .D(n80), .C(Clk), .Q(Dout[14]), .QN(n12) );
  DF3 Dout_reg_13_ ( .D(n81), .C(Clk), .Q(Dout[13]), .QN(n10) );
  DF3 Dout_reg_12_ ( .D(n82), .C(Clk), .Q(Dout[12]), .QN(n8) );
  DF3 Dout_reg_11_ ( .D(n83), .C(Clk), .Q(Dout[11]), .QN(n6) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n58) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n60) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n59) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n84) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n62) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n61) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n87) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n88) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n86) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n85) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n89) );
  DF3 Dout_reg_17_ ( .D(n77), .C(Clk), .Q(Dout[17]), .QN(n18) );
  DF3 Dout_reg_24_ ( .D(n70), .C(Clk), .Q(Dout[24]), .QN(n32) );
  DF3 Dout_reg_18_ ( .D(n76), .C(Clk), .Q(Dout[18]), .QN(n20) );
  DF3 Dout_reg_20_ ( .D(n74), .C(Clk), .Q(Dout[20]), .QN(n24) );
  DF3 Dout_reg_23_ ( .D(n71), .C(Clk), .Q(Dout[23]), .QN(n30) );
  DF3 Dout_reg_22_ ( .D(n72), .C(Clk), .Q(Dout[22]), .QN(n28) );
  DF3 Dout_reg_19_ ( .D(n75), .C(Clk), .Q(Dout[19]), .QN(n22) );
  DF3 Dout_reg_21_ ( .D(n73), .C(Clk), .Q(Dout[21]), .QN(n26) );
  OAI222 U3 ( .A(n85), .B(n360), .C(n362), .D(n394), .Q(n99) );
  OAI222 U4 ( .A(n86), .B(n360), .C(n361), .D(n393), .Q(n98) );
  OAI222 U5 ( .A(n88), .B(n360), .C(n104), .D(n392), .Q(n97) );
  OAI222 U6 ( .A(n87), .B(n360), .C(n362), .D(n391), .Q(n96) );
  OAI222 U7 ( .A(n61), .B(n360), .C(n361), .D(n390), .Q(n95) );
  OAI222 U8 ( .A(n62), .B(n360), .C(n104), .D(n389), .Q(n94) );
  OAI222 U9 ( .A(n84), .B(n360), .C(n362), .D(n388), .Q(n93) );
  OAI222 U10 ( .A(n59), .B(n360), .C(n361), .D(n387), .Q(n92) );
  OAI222 U11 ( .A(n60), .B(n360), .C(n104), .D(n386), .Q(n91) );
  OAI222 U12 ( .A(n58), .B(n360), .C(n362), .D(n385), .Q(n90) );
  OAI222 U13 ( .A(n6), .B(n360), .C(n361), .D(n384), .Q(n83) );
  OAI222 U14 ( .A(n8), .B(n360), .C(n104), .D(n383), .Q(n82) );
  OAI222 U15 ( .A(n10), .B(n360), .C(n362), .D(n382), .Q(n81) );
  OAI222 U16 ( .A(n12), .B(n360), .C(n361), .D(n381), .Q(n80) );
  OAI222 U17 ( .A(n14), .B(n360), .C(n104), .D(n364), .Q(n79) );
  OAI222 U18 ( .A(n16), .B(n360), .C(n362), .D(n366), .Q(n78) );
  OAI222 U19 ( .A(n18), .B(n360), .C(n361), .D(n372), .Q(n77) );
  OAI222 U20 ( .A(n20), .B(n360), .C(n104), .D(n369), .Q(n76) );
  OAI222 U21 ( .A(n22), .B(n360), .C(n362), .D(n367), .Q(n75) );
  OAI222 U22 ( .A(n24), .B(n360), .C(n361), .D(n368), .Q(n74) );
  OAI222 U23 ( .A(n26), .B(n360), .C(n104), .D(n373), .Q(n73) );
  OAI222 U24 ( .A(n28), .B(n360), .C(n362), .D(n370), .Q(n72) );
  OAI222 U25 ( .A(n30), .B(n360), .C(n361), .D(n371), .Q(n71) );
  OAI222 U26 ( .A(n32), .B(n360), .C(n104), .D(n380), .Q(n70) );
  OAI222 U27 ( .A(n35), .B(n360), .C(n362), .D(n374), .Q(n69) );
  OAI222 U28 ( .A(n47), .B(n360), .C(n361), .D(n375), .Q(n68) );
  OAI222 U29 ( .A(n49), .B(n360), .C(n104), .D(n379), .Q(n67) );
  OAI222 U30 ( .A(n51), .B(n360), .C(n362), .D(n376), .Q(n66) );
  OAI222 U31 ( .A(n53), .B(n360), .C(n361), .D(n365), .Q(n65) );
  OAI222 U32 ( .A(n55), .B(n360), .C(n104), .D(n378), .Q(n64) );
  OAI222 U33 ( .A(n57), .B(n360), .C(n377), .D(n362), .Q(n63) );
  OAI222 U34 ( .A(n89), .B(n360), .C(n361), .D(n395), .Q(n100) );
  DF1 Dout_reg_28_ ( .D(n66), .C(Clk), .Q(Dout[28]), .QN(n51) );
  DF1 Dout_reg_25_ ( .D(n69), .C(Clk), .Q(Dout[25]), .QN(n35) );
  DF1 Dout_reg_31_ ( .D(n63), .C(Clk), .Q(Dout[31]), .QN(n57) );
  DF1 Dout_reg_30_ ( .D(n64), .C(Clk), .Q(Dout[30]), .QN(n55) );
  DF3 Dout_reg_27_ ( .D(n67), .C(Clk), .Q(Dout[27]), .QN(n49) );
  DF3 Dout_reg_26_ ( .D(n68), .C(Clk), .Q(Dout[26]), .QN(n47) );
  DF1 Dout_reg_29_ ( .D(n65), .C(Clk), .Q(Dout[29]), .QN(n53) );
  INV4 U35 ( .A(Din[27]), .Q(n379) );
  INV3 U36 ( .A(Din[17]), .Q(n372) );
  INV3 U37 ( .A(Din[28]), .Q(n376) );
  INV3 U38 ( .A(Din[20]), .Q(n368) );
  INV3 U39 ( .A(Din[21]), .Q(n373) );
  INV3 U40 ( .A(Din[29]), .Q(n365) );
  INV4 U41 ( .A(Din[31]), .Q(n377) );
  INV3 U42 ( .A(Din[30]), .Q(n378) );
  CLKIN2 U43 ( .A(Din[8]), .Q(n387) );
  INV3 U44 ( .A(Din[12]), .Q(n383) );
  INV3 U45 ( .A(Din[10]), .Q(n385) );
  INV3 U46 ( .A(Din[11]), .Q(n384) );
  INV3 U47 ( .A(Din[9]), .Q(n386) );
  INV2 U48 ( .A(Din[25]), .Q(n374) );
  INV2 U49 ( .A(Din[26]), .Q(n375) );
  INV2 U50 ( .A(Din[23]), .Q(n371) );
  INV2 U51 ( .A(Din[19]), .Q(n367) );
  INV2 U52 ( .A(Din[22]), .Q(n370) );
  INV2 U53 ( .A(Din[16]), .Q(n366) );
  INV2 U54 ( .A(Din[24]), .Q(n380) );
  INV2 U55 ( .A(Din[18]), .Q(n369) );
  INV2 U56 ( .A(Din[14]), .Q(n381) );
  INV2 U57 ( .A(Din[13]), .Q(n382) );
  INV2 U58 ( .A(Din[15]), .Q(n364) );
  INV2 U59 ( .A(Din[6]), .Q(n389) );
  NAND22 U60 ( .A(n363), .B(n360), .Q(n361) );
  NAND22 U61 ( .A(n363), .B(n360), .Q(n362) );
  NAND22 U62 ( .A(n363), .B(n360), .Q(n104) );
  INV3 U63 ( .A(Reset), .Q(n363) );
  INV3 U64 ( .A(n105), .Q(n360) );
  INV3 U65 ( .A(Din[7]), .Q(n388) );
  INV3 U66 ( .A(Din[2]), .Q(n393) );
  INV3 U67 ( .A(Din[4]), .Q(n391) );
  INV3 U68 ( .A(Din[5]), .Q(n390) );
  INV3 U69 ( .A(Din[1]), .Q(n394) );
  INV3 U70 ( .A(Din[3]), .Q(n392) );
  INV3 U71 ( .A(Din[0]), .Q(n395) );
  NOR21 U72 ( .A(Load), .B(Reset), .Q(n105) );
endmodule


module adder_9_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n198, n203, n204, n205, n206, n207, n208, n209, n212, n213,
         n214, n219, n220, n221, n222, n223, n224, n225, n226, n227, n230,
         n231, n232, n239, n240, n242, n243, n245, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n265, n266, n268, n269, n270, n271, n272, n273, n274, n275,
         n277, n278, n279, n280, n281, n423, n426, n429, n430, n500, n501,
         n505, n506, n507, n508, n509, n510, n513, n585, n588, n589, n590,
         n595, n596, n597, n677, n759, n760, n761, n764, n765, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934;

  OAI212 U77 ( .A(n91), .B(n853), .C(n92), .Q(n90) );
  OAI212 U91 ( .A(n102), .B(n853), .C(n103), .Q(n101) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n853), .C(n121), .Q(n119) );
  OAI212 U141 ( .A(n140), .B(n853), .C(n141), .Q(n139) );
  OAI212 U165 ( .A(n158), .B(n853), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n856), .B(n853), .C(n862), .Q(n164) );
  AOI212 U195 ( .A(n507), .B(n179), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U219 ( .A(n870), .B(n888), .C(n198), .Q(n196) );
  OAI212 U233 ( .A(n208), .B(n888), .C(n209), .Q(n207) );
  OAI212 U257 ( .A(n226), .B(n888), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n884), .B(n888), .C(n882), .Q(n232) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  AOI212 U389 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U417 ( .A(n64), .B(n853), .C(n65), .Q(n63) );
  OAI212 U427 ( .A(n129), .B(n853), .C(n130), .Q(n128) );
  OAI212 U463 ( .A(n176), .B(n853), .C(n177), .Q(n175) );
  AOI212 U390 ( .A(n509), .B(n760), .C(n590), .Q(n510) );
  OAI212 U399 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U400 ( .A(n274), .B(n898), .C(n275), .Q(n273) );
  OAI212 U501 ( .A(n188), .B(n888), .C(n189), .Q(n187) );
  OAI212 U495 ( .A(n858), .B(n853), .C(n864), .Q(n108) );
  OAI212 U535 ( .A(n145), .B(n920), .C(n138), .Q(n136) );
  OAI212 U664 ( .A(n886), .B(n888), .C(n245), .Q(n243) );
  AOI212 U388 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U446 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U404 ( .A(n42), .B(n853), .C(n43), .Q(n41) );
  OAI212 U401 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U406 ( .A(n245), .B(n513), .C(n242), .Q(n509) );
  OAI212 U437 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U449 ( .A(n53), .B(n853), .C(n54), .Q(n52) );
  OAI212 U476 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U482 ( .A(n73), .B(n853), .C(n74), .Q(n72) );
  XNR22 U494 ( .A(n23), .B(n187), .Q(SUM[15]) );
  XNR22 U497 ( .A(n27), .B(n225), .Q(SUM[11]) );
  OAI212 U498 ( .A(n82), .B(n853), .C(n83), .Q(n81) );
  XNR22 U503 ( .A(n28), .B(n232), .Q(SUM[10]) );
  XOR22 U505 ( .A(n22), .B(n853), .Q(SUM[16]) );
  OAI212 U508 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  XNR22 U518 ( .A(n25), .B(n207), .Q(SUM[13]) );
  XNR22 U533 ( .A(n24), .B(n196), .Q(SUM[14]) );
  OAI212 U439 ( .A(n126), .B(n915), .C(n127), .Q(n123) );
  OAI212 U483 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U527 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  INV3 U349 ( .A(n423), .Q(n870) );
  CLKIN4 U350 ( .A(A[8]), .Q(n933) );
  NAND23 U351 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND28 U352 ( .A(n585), .B(n174), .Q(n172) );
  XNR22 U353 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NOR24 U354 ( .A(n252), .B(n255), .Q(n250) );
  INV1 U355 ( .A(n255), .Q(n890) );
  OAI211 U356 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NAND24 U357 ( .A(n500), .B(n501), .Q(SUM[9]) );
  CLKIN6 U358 ( .A(n157), .Q(n860) );
  NAND22 U359 ( .A(n157), .B(n19), .Q(n595) );
  AOI212 U360 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NOR24 U361 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NAND26 U362 ( .A(n764), .B(n765), .Q(SUM[18]) );
  NOR22 U363 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR24 U364 ( .A(n212), .B(n205), .Q(n203) );
  INV1 U365 ( .A(n194), .Q(n867) );
  NOR22 U366 ( .A(n194), .B(n871), .Q(n190) );
  NOR24 U367 ( .A(n185), .B(n194), .Q(n183) );
  NOR23 U368 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND23 U369 ( .A(n171), .B(n153), .Q(n151) );
  NOR22 U370 ( .A(n155), .B(n162), .Q(n153) );
  NAND22 U371 ( .A(n875), .B(n224), .Q(n27) );
  NOR22 U372 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NOR22 U373 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NAND24 U374 ( .A(n203), .B(n183), .Q(n761) );
  INV6 U375 ( .A(n759), .Q(n886) );
  INV3 U376 ( .A(n243), .Q(n885) );
  NOR22 U377 ( .A(n761), .B(n219), .Q(n179) );
  NOR23 U378 ( .A(n79), .B(n88), .Q(n77) );
  NOR21 U379 ( .A(n70), .B(n6), .Q(n66) );
  INV3 U380 ( .A(n175), .Q(n861) );
  NOR22 U381 ( .A(n920), .B(n144), .Q(n135) );
  BUF6 U382 ( .A(n213), .Q(n849) );
  NAND24 U383 ( .A(n239), .B(n221), .Q(n219) );
  NOR22 U384 ( .A(n99), .B(n106), .Q(n97) );
  INV3 U385 ( .A(n151), .Q(n857) );
  NAND22 U386 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND24 U387 ( .A(n887), .B(n933), .Q(n759) );
  NOR23 U391 ( .A(B[15]), .B(A[15]), .Q(n185) );
  INV3 U392 ( .A(n90), .Q(n859) );
  NAND22 U393 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND22 U394 ( .A(A[11]), .B(B[11]), .Q(n224) );
  CLKIN1 U395 ( .A(n136), .Q(n915) );
  AOI211 U396 ( .A(n876), .B(n203), .C(n426), .Q(n198) );
  NAND21 U397 ( .A(n924), .B(n100), .Q(n13) );
  CLKIN2 U398 ( .A(n230), .Q(n880) );
  OAI210 U402 ( .A(n194), .B(n868), .C(n195), .Q(n191) );
  NAND22 U403 ( .A(n26), .B(n214), .Q(n505) );
  NAND26 U405 ( .A(n429), .B(n430), .Q(SUM[17]) );
  NOR23 U407 ( .A(B[11]), .B(A[11]), .Q(n597) );
  NOR23 U408 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND22 U409 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND20 U410 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NOR21 U411 ( .A(n88), .B(n904), .Q(n84) );
  OAI211 U412 ( .A(n205), .B(n849), .C(n206), .Q(n426) );
  AOI212 U413 ( .A(n851), .B(n97), .C(n98), .Q(n92) );
  NAND21 U414 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND24 U415 ( .A(n505), .B(n506), .Q(SUM[12]) );
  NAND21 U416 ( .A(A[21]), .B(B[21]), .Q(n138) );
  INV6 U418 ( .A(n848), .Q(n902) );
  AOI211 U419 ( .A(n172), .B(n911), .C(n909), .Q(n159) );
  NAND21 U420 ( .A(n20), .B(n164), .Q(n764) );
  NAND21 U421 ( .A(A[15]), .B(B[15]), .Q(n186) );
  AOI211 U422 ( .A(n863), .B(n122), .C(n123), .Q(n121) );
  NAND22 U423 ( .A(n857), .B(n122), .Q(n120) );
  INV3 U424 ( .A(n152), .Q(n863) );
  NAND28 U425 ( .A(n595), .B(n596), .Q(SUM[19]) );
  NOR22 U426 ( .A(n597), .B(n230), .Q(n760) );
  OAI211 U428 ( .A(n231), .B(n223), .C(n224), .Q(n590) );
  NAND24 U429 ( .A(n865), .B(n902), .Q(n585) );
  NAND20 U430 ( .A(A[25]), .B(B[25]), .Q(n100) );
  INV1 U431 ( .A(n212), .Q(n874) );
  NAND24 U432 ( .A(n910), .B(n855), .Q(n765) );
  CLKIN4 U433 ( .A(n164), .Q(n855) );
  NAND21 U434 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND21 U435 ( .A(n12), .B(n90), .Q(n588) );
  NAND22 U436 ( .A(A[17]), .B(B[17]), .Q(n174) );
  INV3 U438 ( .A(n106), .Q(n903) );
  NOR23 U440 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND21 U441 ( .A(A[26]), .B(B[26]), .Q(n89) );
  OAI212 U442 ( .A(n245), .B(n513), .C(n242), .Q(n240) );
  NOR24 U443 ( .A(B[9]), .B(A[9]), .Q(n513) );
  AOI212 U444 ( .A(n851), .B(n903), .C(n906), .Q(n103) );
  NAND26 U445 ( .A(n860), .B(n918), .Q(n596) );
  NAND26 U447 ( .A(n861), .B(n901), .Q(n430) );
  INV6 U448 ( .A(n850), .Q(n851) );
  NAND21 U450 ( .A(n919), .B(n156), .Q(n19) );
  NAND22 U451 ( .A(n258), .B(n250), .Q(n248) );
  NOR24 U452 ( .A(B[7]), .B(A[7]), .Q(n252) );
  OAI211 U453 ( .A(n219), .B(n888), .C(n510), .Q(n214) );
  CLKIN3 U454 ( .A(n219), .Q(n878) );
  INV6 U455 ( .A(n112), .Q(n850) );
  CLKIN6 U456 ( .A(n850), .Q(n852) );
  NAND22 U457 ( .A(n111), .B(n84), .Q(n82) );
  OAI212 U458 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI211 U459 ( .A(n248), .B(n268), .C(n249), .Q(n507) );
  OAI211 U460 ( .A(n88), .B(n907), .C(n89), .Q(n85) );
  INV2 U461 ( .A(n98), .Q(n907) );
  NAND22 U462 ( .A(n203), .B(n183), .Q(n181) );
  NAND23 U464 ( .A(n921), .B(n934), .Q(n677) );
  INV2 U465 ( .A(A[21]), .Q(n934) );
  AOI211 U466 ( .A(n863), .B(n135), .C(n136), .Q(n130) );
  AOI211 U467 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  XNR22 U468 ( .A(n8), .B(n52), .Q(SUM[30]) );
  OAI211 U469 ( .A(n205), .B(n849), .C(n206), .Q(n204) );
  NOR22 U470 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NAND21 U471 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NOR24 U472 ( .A(n113), .B(n151), .Q(n111) );
  NAND24 U473 ( .A(n135), .B(n115), .Q(n113) );
  NAND20 U474 ( .A(n677), .B(n138), .Q(n17) );
  NOR22 U475 ( .A(n597), .B(n230), .Q(n221) );
  NAND22 U477 ( .A(n175), .B(n21), .Q(n429) );
  INV6 U478 ( .A(n677), .Q(n920) );
  OAI212 U479 ( .A(n151), .B(n853), .C(n847), .Q(n146) );
  NOR22 U480 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND24 U481 ( .A(n97), .B(n77), .Q(n6) );
  INV2 U484 ( .A(n863), .Q(n847) );
  NAND24 U485 ( .A(n588), .B(n589), .Q(SUM[26]) );
  NOR22 U486 ( .A(n117), .B(n126), .Q(n115) );
  NOR20 U487 ( .A(n219), .B(n871), .Q(n423) );
  CLKIN3 U488 ( .A(n203), .Q(n871) );
  AOI211 U489 ( .A(n876), .B(n190), .C(n191), .Q(n189) );
  NAND21 U490 ( .A(n869), .B(n206), .Q(n25) );
  NAND21 U491 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND22 U492 ( .A(n903), .B(n107), .Q(n14) );
  NAND21 U493 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NOR22 U496 ( .A(B[17]), .B(A[17]), .Q(n173) );
  INV0 U499 ( .A(n117), .Q(n916) );
  CLKIN2 U500 ( .A(n135), .Q(n913) );
  AOI211 U502 ( .A(n852), .B(n55), .C(n56), .Q(n54) );
  XNR22 U504 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND22 U506 ( .A(n911), .B(n163), .Q(n20) );
  NAND22 U507 ( .A(A[18]), .B(B[18]), .Q(n163) );
  OAI211 U509 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NAND22 U510 ( .A(n111), .B(n97), .Q(n91) );
  CLKIN3 U511 ( .A(n111), .Q(n858) );
  NAND22 U512 ( .A(n111), .B(n66), .Q(n64) );
  XNR22 U513 ( .A(n16), .B(n128), .Q(SUM[22]) );
  XNR22 U514 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U515 ( .A(n9), .B(n63), .Q(SUM[29]) );
  INV3 U516 ( .A(n70), .Q(n931) );
  OAI211 U517 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  NOR22 U519 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NAND22 U520 ( .A(n111), .B(n55), .Q(n53) );
  NOR21 U521 ( .A(n930), .B(n6), .Q(n55) );
  XNR22 U522 ( .A(n10), .B(n72), .Q(SUM[28]) );
  NOR21 U523 ( .A(n61), .B(n70), .Q(n59) );
  NOR22 U524 ( .A(B[29]), .B(A[29]), .Q(n61) );
  XNR22 U525 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U526 ( .A(n15), .B(n119), .Q(SUM[23]) );
  XNR22 U528 ( .A(n13), .B(n101), .Q(SUM[25]) );
  BUF6 U529 ( .A(n173), .Q(n848) );
  NAND20 U530 ( .A(n239), .B(n880), .Q(n226) );
  CLKIN0 U531 ( .A(n239), .Q(n884) );
  NOR24 U532 ( .A(n513), .B(n886), .Q(n239) );
  NAND21 U534 ( .A(n857), .B(n135), .Q(n129) );
  AOI210 U536 ( .A(n895), .B(n258), .C(n259), .Q(n257) );
  INV2 U537 ( .A(n5), .Q(n908) );
  INV1 U538 ( .A(n6), .Q(n905) );
  CLKIN3 U539 ( .A(B[21]), .Q(n921) );
  CLKIN3 U540 ( .A(B[8]), .Q(n887) );
  NAND21 U541 ( .A(n111), .B(n903), .Q(n102) );
  NAND21 U542 ( .A(n878), .B(n190), .Q(n188) );
  AOI211 U543 ( .A(n852), .B(n66), .C(n67), .Q(n65) );
  NAND20 U544 ( .A(n866), .B(n186), .Q(n23) );
  INV0 U545 ( .A(n163), .Q(n909) );
  CLKIN12 U546 ( .A(n247), .Q(n888) );
  NAND21 U547 ( .A(n29), .B(n243), .Q(n500) );
  INV2 U548 ( .A(n29), .Q(n881) );
  CLKIN3 U549 ( .A(n59), .Q(n930) );
  AOI212 U550 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  AOI211 U551 ( .A(n876), .B(n874), .C(n872), .Q(n209) );
  INV2 U552 ( .A(n97), .Q(n904) );
  NAND20 U553 ( .A(n854), .B(n177), .Q(n22) );
  AOI212 U554 ( .A(n760), .B(n240), .C(n222), .Q(n220) );
  INV0 U555 ( .A(n205), .Q(n869) );
  NOR22 U556 ( .A(n848), .B(n176), .Q(n171) );
  INV0 U557 ( .A(n126), .Q(n917) );
  CLKIN0 U558 ( .A(n162), .Q(n911) );
  NAND20 U559 ( .A(n923), .B(n89), .Q(n12) );
  INV0 U560 ( .A(n88), .Q(n923) );
  INV2 U561 ( .A(n271), .Q(n894) );
  NAND20 U562 ( .A(n867), .B(n195), .Q(n24) );
  NAND20 U563 ( .A(n902), .B(n174), .Q(n21) );
  INV0 U564 ( .A(n185), .Q(n866) );
  NAND21 U565 ( .A(n874), .B(n849), .Q(n26) );
  INV2 U566 ( .A(n265), .Q(n893) );
  INV2 U567 ( .A(n274), .Q(n896) );
  INV2 U568 ( .A(n260), .Q(n891) );
  OAI210 U569 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  NOR20 U570 ( .A(n271), .B(n274), .Q(n269) );
  NAND20 U571 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U572 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND20 U573 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U574 ( .A(n111), .B(n905), .Q(n73) );
  NAND20 U575 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U576 ( .A(n214), .Q(n877) );
  INV3 U577 ( .A(n852), .Q(n864) );
  INV3 U578 ( .A(n172), .Q(n862) );
  INV3 U579 ( .A(n171), .Q(n856) );
  INV3 U580 ( .A(n60), .Q(n929) );
  NOR20 U581 ( .A(n46), .B(n6), .Q(n44) );
  NAND22 U582 ( .A(n922), .B(n859), .Q(n589) );
  INV3 U583 ( .A(n12), .Q(n922) );
  AOI211 U584 ( .A(n852), .B(n905), .C(n908), .Q(n74) );
  INV3 U585 ( .A(n21), .Q(n901) );
  NAND22 U586 ( .A(n873), .B(n877), .Q(n506) );
  INV3 U587 ( .A(n26), .Q(n873) );
  INV3 U588 ( .A(n20), .Q(n910) );
  NAND22 U589 ( .A(n881), .B(n885), .Q(n501) );
  INV3 U590 ( .A(n19), .Q(n918) );
  NAND22 U591 ( .A(n878), .B(n874), .Q(n208) );
  INV3 U592 ( .A(n510), .Q(n876) );
  CLKIN0 U593 ( .A(n509), .Q(n882) );
  INV3 U594 ( .A(n268), .Q(n895) );
  INV3 U595 ( .A(n277), .Q(n898) );
  NAND22 U596 ( .A(n171), .B(n911), .Q(n158) );
  XOR21 U597 ( .A(n30), .B(n888), .Q(SUM[8]) );
  NAND20 U598 ( .A(n759), .B(n245), .Q(n30) );
  XOR21 U599 ( .A(n32), .B(n508), .Q(SUM[6]) );
  NAND20 U600 ( .A(n890), .B(n256), .Q(n32) );
  AOI210 U601 ( .A(n895), .B(n258), .C(n259), .Q(n508) );
  XOR21 U602 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U603 ( .A(n895), .B(n893), .C(n892), .Q(n262) );
  NAND22 U604 ( .A(n891), .B(n261), .Q(n33) );
  INV3 U605 ( .A(n266), .Q(n892) );
  XOR21 U606 ( .A(n36), .B(n898), .Q(SUM[2]) );
  NAND22 U607 ( .A(n896), .B(n275), .Q(n36) );
  XNR21 U608 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U609 ( .A(n889), .B(n253), .Q(n31) );
  INV0 U610 ( .A(n252), .Q(n889) );
  NAND20 U611 ( .A(n931), .B(n71), .Q(n10) );
  NAND22 U612 ( .A(n932), .B(n80), .Q(n11) );
  INV3 U613 ( .A(n79), .Q(n932) );
  NAND22 U614 ( .A(n928), .B(n62), .Q(n9) );
  INV3 U615 ( .A(n61), .Q(n928) );
  NAND22 U616 ( .A(n926), .B(n51), .Q(n8) );
  XNR21 U617 ( .A(n34), .B(n895), .Q(SUM[4]) );
  NAND22 U618 ( .A(n893), .B(n266), .Q(n34) );
  XNR21 U619 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U620 ( .A(n894), .B(n272), .Q(n35) );
  XOR21 U621 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U622 ( .A(n897), .B(n279), .Q(n37) );
  INV3 U623 ( .A(n278), .Q(n897) );
  NAND20 U624 ( .A(n880), .B(n231), .Q(n28) );
  INV3 U625 ( .A(n176), .Q(n854) );
  NAND20 U626 ( .A(n912), .B(n145), .Q(n18) );
  NAND20 U627 ( .A(n917), .B(n127), .Q(n16) );
  INV0 U628 ( .A(n223), .Q(n875) );
  AOI210 U629 ( .A(n60), .B(n926), .C(n927), .Q(n47) );
  INV3 U630 ( .A(n51), .Q(n927) );
  INV0 U631 ( .A(n99), .Q(n924) );
  NAND22 U632 ( .A(n857), .B(n912), .Q(n140) );
  NOR21 U633 ( .A(n126), .B(n913), .Q(n122) );
  NAND22 U634 ( .A(n916), .B(n118), .Q(n15) );
  INV3 U635 ( .A(n107), .Q(n906) );
  INV3 U636 ( .A(n155), .Q(n919) );
  CLKIN3 U637 ( .A(n177), .Q(n865) );
  NAND21 U638 ( .A(n883), .B(n242), .Q(n29) );
  INV0 U639 ( .A(n513), .Q(n883) );
  AOI210 U640 ( .A(n509), .B(n880), .C(n879), .Q(n227) );
  INV0 U641 ( .A(n231), .Q(n879) );
  AOI211 U642 ( .A(n863), .B(n912), .C(n914), .Q(n141) );
  INV0 U643 ( .A(n145), .Q(n914) );
  INV3 U644 ( .A(n426), .Q(n868) );
  INV3 U645 ( .A(n849), .Q(n872) );
  NAND20 U646 ( .A(n59), .B(n926), .Q(n46) );
  AOI211 U647 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR20 U648 ( .A(n260), .B(n265), .Q(n258) );
  XNR21 U649 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U650 ( .A(n925), .B(n40), .Q(n7) );
  NAND20 U651 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR21 U652 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR21 U653 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR20 U654 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR20 U655 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR20 U656 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR20 U657 ( .A(B[1]), .B(A[1]), .Q(n278) );
  INV3 U658 ( .A(n38), .Q(SUM[0]) );
  NAND22 U659 ( .A(n900), .B(n281), .Q(n38) );
  INV3 U660 ( .A(n280), .Q(n900) );
  NOR20 U661 ( .A(B[0]), .B(A[0]), .Q(n280) );
  INV3 U662 ( .A(n39), .Q(n925) );
  INV3 U663 ( .A(n50), .Q(n926) );
  NOR20 U665 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND20 U666 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U667 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U668 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U669 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND21 U670 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND21 U671 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND22 U672 ( .A(A[7]), .B(B[7]), .Q(n253) );
  OAI210 U673 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI210 U674 ( .A(n930), .B(n5), .C(n929), .Q(n56) );
  INV3 U675 ( .A(n144), .Q(n912) );
  AOI211 U676 ( .A(n851), .B(n84), .C(n85), .Q(n83) );
  NOR21 U677 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND22 U678 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NOR22 U679 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR21 U680 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND22 U681 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND22 U682 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NOR22 U683 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR21 U684 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND22 U685 ( .A(A[16]), .B(B[16]), .Q(n177) );
  AOI210 U686 ( .A(n852), .B(n44), .C(n45), .Q(n43) );
  NOR21 U687 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR22 U688 ( .A(B[11]), .B(A[11]), .Q(n223) );
  BUF15 U689 ( .A(n178), .Q(n853) );
endmodule


module adder_9 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_9_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_8_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n85, n88, n89, n90, n91, n92, n98, n99, n100, n101, n102, n103, n106,
         n107, n108, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n126, n127, n128, n129, n130, n135, n136,
         n138, n139, n140, n141, n144, n145, n146, n151, n153, n154, n155,
         n156, n157, n158, n159, n162, n163, n164, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n194, n195, n196, n197, n198,
         n203, n204, n205, n206, n207, n208, n209, n212, n213, n214, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n230, n231, n232,
         n239, n240, n241, n242, n243, n244, n245, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n265, n266, n268, n269, n270, n271, n272, n273, n274, n275,
         n277, n278, n279, n280, n281, n418, n426, n428, n501, n508, n511,
         n515, n580, n584, n588, n592, n661, n674, n745, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n898;

  OAI212 U105 ( .A(n508), .B(n113), .C(n114), .Q(n112) );
  OAI212 U201 ( .A(n185), .B(n195), .C(n186), .Q(n184) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U292 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n896), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U380 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  AOI212 U492 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U456 ( .A(n418), .B(n865), .C(n866), .Q(n56) );
  OAI212 U510 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U413 ( .A(n830), .B(n102), .C(n103), .Q(n101) );
  OAI212 U454 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  OAI212 U480 ( .A(n661), .B(n145), .C(n138), .Q(n136) );
  OAI212 U519 ( .A(n173), .B(n177), .C(n174), .Q(n172) );
  OAI212 U526 ( .A(n79), .B(n89), .C(n80), .Q(n78) );
  AOI212 U546 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  AOI212 U549 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI212 U353 ( .A(n129), .B(n830), .C(n130), .Q(n128) );
  OAI212 U496 ( .A(n850), .B(n830), .C(n847), .Q(n164) );
  OAI212 U497 ( .A(n158), .B(n830), .C(n159), .Q(n157) );
  OAI212 U502 ( .A(n830), .B(n73), .C(n74), .Q(n72) );
  NOR24 U516 ( .A(n822), .B(n144), .Q(n135) );
  OAI212 U499 ( .A(n188), .B(n887), .C(n189), .Q(n187) );
  OAI212 U500 ( .A(n226), .B(n887), .C(n227), .Q(n225) );
  OAI212 U501 ( .A(n883), .B(n887), .C(n884), .Q(n232) );
  BUF2 U349 ( .A(n185), .Q(n816) );
  NOR24 U350 ( .A(A[12]), .B(B[12]), .Q(n212) );
  BUF2 U351 ( .A(n127), .Q(n823) );
  NOR23 U352 ( .A(n223), .B(n230), .Q(n221) );
  NOR23 U354 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR23 U355 ( .A(A[27]), .B(B[27]), .Q(n79) );
  NAND28 U356 ( .A(n588), .B(n100), .Q(n98) );
  INV1 U357 ( .A(n220), .Q(n877) );
  INV2 U358 ( .A(n6), .Q(n840) );
  NOR24 U359 ( .A(n70), .B(n6), .Q(n66) );
  INV2 U360 ( .A(n508), .Q(n848) );
  INV0 U361 ( .A(n816), .Q(n832) );
  NAND23 U362 ( .A(B[16]), .B(A[16]), .Q(n177) );
  NAND23 U363 ( .A(n171), .B(n153), .Q(n151) );
  NOR23 U364 ( .A(n155), .B(n162), .Q(n153) );
  NAND22 U365 ( .A(B[13]), .B(A[13]), .Q(n206) );
  NAND22 U366 ( .A(n851), .B(n862), .Q(n140) );
  NOR24 U367 ( .A(n185), .B(n194), .Q(n183) );
  NOR24 U368 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR23 U369 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR23 U370 ( .A(n828), .B(n78), .Q(n418) );
  NAND24 U371 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NOR24 U372 ( .A(n212), .B(n817), .Q(n203) );
  NOR24 U373 ( .A(B[13]), .B(A[13]), .Q(n817) );
  NAND22 U374 ( .A(n818), .B(n819), .Q(n821) );
  NAND24 U375 ( .A(n511), .B(n71), .Q(n67) );
  NOR23 U376 ( .A(n181), .B(n219), .Q(n179) );
  INV3 U377 ( .A(n107), .Q(n867) );
  NOR23 U378 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR22 U379 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR23 U381 ( .A(A[18]), .B(B[18]), .Q(n162) );
  NOR22 U382 ( .A(n173), .B(n176), .Q(n171) );
  NOR23 U383 ( .A(A[11]), .B(B[11]), .Q(n223) );
  NAND24 U384 ( .A(n203), .B(n183), .Q(n181) );
  NAND23 U385 ( .A(n842), .B(n831), .Q(n592) );
  INV3 U386 ( .A(n418), .Q(n836) );
  NAND22 U387 ( .A(n580), .B(n823), .Q(n123) );
  NAND22 U388 ( .A(B[18]), .B(A[18]), .Q(n163) );
  AOI211 U389 ( .A(n877), .B(n875), .C(n876), .Q(n209) );
  NAND22 U390 ( .A(n820), .B(n821), .Q(SUM[17]) );
  NOR23 U391 ( .A(A[21]), .B(B[21]), .Q(n822) );
  NOR23 U392 ( .A(A[21]), .B(B[21]), .Q(n661) );
  NAND22 U393 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U394 ( .A(n846), .B(n80), .Q(n11) );
  NAND21 U395 ( .A(n21), .B(n175), .Q(n820) );
  INV0 U396 ( .A(n21), .Q(n818) );
  INV3 U397 ( .A(n175), .Q(n819) );
  INV6 U398 ( .A(n77), .Q(n839) );
  AOI212 U399 ( .A(n60), .B(n833), .C(n834), .Q(n47) );
  NAND22 U400 ( .A(n833), .B(n51), .Q(n8) );
  NOR24 U401 ( .A(A[15]), .B(B[15]), .Q(n185) );
  NOR23 U402 ( .A(B[28]), .B(A[28]), .Q(n70) );
  AOI211 U403 ( .A(n829), .B(n840), .C(n836), .Q(n74) );
  INV8 U404 ( .A(n829), .Q(n843) );
  NAND22 U405 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR21 U406 ( .A(n194), .B(n874), .Q(n190) );
  INV1 U407 ( .A(n194), .Q(n871) );
  OAI210 U408 ( .A(n194), .B(n872), .C(n195), .Q(n191) );
  NAND22 U409 ( .A(B[19]), .B(A[19]), .Q(n156) );
  NAND24 U410 ( .A(n854), .B(n868), .Q(n501) );
  INV0 U411 ( .A(n204), .Q(n872) );
  OAI211 U412 ( .A(n145), .B(n661), .C(n138), .Q(n426) );
  AOI211 U414 ( .A(n848), .B(n122), .C(n123), .Q(n121) );
  NOR24 U415 ( .A(B[24]), .B(A[24]), .Q(n106) );
  INV4 U416 ( .A(n98), .Q(n827) );
  INV8 U417 ( .A(n501), .Q(n853) );
  INV6 U418 ( .A(n98), .Q(n852) );
  INV4 U419 ( .A(n5), .Q(n835) );
  XNR22 U420 ( .A(n13), .B(n101), .Q(SUM[25]) );
  NAND22 U421 ( .A(B[17]), .B(A[17]), .Q(n174) );
  NOR23 U422 ( .A(n151), .B(n113), .Q(n111) );
  CLKIN2 U423 ( .A(n126), .Q(n844) );
  NOR22 U424 ( .A(A[8]), .B(B[8]), .Q(n244) );
  NOR23 U425 ( .A(n46), .B(n6), .Q(n44) );
  CLKIN6 U426 ( .A(n50), .Q(n833) );
  NOR22 U427 ( .A(B[30]), .B(A[30]), .Q(n50) );
  OAI211 U428 ( .A(n219), .B(n887), .C(n220), .Q(n214) );
  INV6 U429 ( .A(n106), .Q(n868) );
  NOR24 U430 ( .A(n839), .B(n852), .Q(n515) );
  CLKIN3 U431 ( .A(n66), .Q(n841) );
  INV1 U432 ( .A(n144), .Q(n862) );
  NAND22 U433 ( .A(n838), .B(n853), .Q(n584) );
  INV4 U434 ( .A(n584), .Q(n837) );
  INV0 U435 ( .A(n173), .Q(n860) );
  OAI210 U436 ( .A(n177), .B(n173), .C(n174), .Q(n428) );
  XNR22 U437 ( .A(n10), .B(n72), .Q(SUM[28]) );
  INV0 U438 ( .A(n155), .Q(n857) );
  NOR24 U439 ( .A(n827), .B(n839), .Q(n828) );
  NAND22 U440 ( .A(n111), .B(n837), .Q(n82) );
  CLKIN3 U441 ( .A(n247), .Q(n887) );
  OAI211 U442 ( .A(n197), .B(n887), .C(n198), .Q(n196) );
  OAI211 U443 ( .A(n208), .B(n887), .C(n209), .Q(n207) );
  NAND21 U444 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND24 U445 ( .A(n59), .B(n833), .Q(n46) );
  OAI212 U446 ( .A(n845), .B(n830), .C(n843), .Q(n108) );
  NAND21 U447 ( .A(n851), .B(n122), .Q(n120) );
  AOI212 U448 ( .A(n829), .B(n44), .C(n45), .Q(n43) );
  NAND20 U449 ( .A(n869), .B(n71), .Q(n10) );
  NAND22 U450 ( .A(A[28]), .B(B[28]), .Q(n71) );
  INV3 U451 ( .A(n60), .Q(n866) );
  NAND23 U452 ( .A(n835), .B(n869), .Q(n511) );
  NAND22 U453 ( .A(n111), .B(n66), .Q(n64) );
  INV3 U455 ( .A(n64), .Q(n842) );
  NAND21 U457 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NOR24 U458 ( .A(n67), .B(n674), .Q(n65) );
  NOR23 U459 ( .A(A[23]), .B(B[23]), .Q(n117) );
  NOR23 U460 ( .A(A[23]), .B(B[23]), .Q(n745) );
  INV0 U461 ( .A(n79), .Q(n846) );
  OAI212 U462 ( .A(n830), .B(n120), .C(n121), .Q(n119) );
  NAND22 U463 ( .A(n111), .B(n44), .Q(n42) );
  OAI210 U464 ( .A(n88), .B(n852), .C(n89), .Q(n85) );
  CLKIN3 U465 ( .A(n88), .Q(n838) );
  CLKBU15 U466 ( .A(n178), .Q(n830) );
  NOR24 U467 ( .A(n865), .B(n6), .Q(n55) );
  XNR22 U468 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI212 U469 ( .A(n830), .B(n91), .C(n92), .Q(n90) );
  NAND21 U470 ( .A(B[27]), .B(A[27]), .Q(n80) );
  NOR24 U471 ( .A(n78), .B(n515), .Q(n5) );
  NAND24 U472 ( .A(n867), .B(n854), .Q(n588) );
  NAND24 U473 ( .A(n824), .B(n825), .Q(n826) );
  OAI211 U474 ( .A(n176), .B(n830), .C(n177), .Q(n175) );
  NOR24 U475 ( .A(n843), .B(n841), .Q(n674) );
  NOR22 U476 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND24 U477 ( .A(n239), .B(n221), .Q(n219) );
  NOR22 U478 ( .A(n241), .B(n244), .Q(n239) );
  INV6 U479 ( .A(n99), .Q(n854) );
  AOI210 U481 ( .A(n848), .B(n135), .C(n426), .Q(n130) );
  NAND21 U482 ( .A(n851), .B(n135), .Q(n129) );
  INV3 U483 ( .A(n135), .Q(n856) );
  OAI212 U484 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U485 ( .A(n244), .B(n887), .C(n245), .Q(n243) );
  INV0 U486 ( .A(n822), .Q(n855) );
  AOI212 U487 ( .A(n829), .B(n55), .C(n56), .Q(n54) );
  NOR24 U488 ( .A(n745), .B(n126), .Q(n115) );
  INV1 U489 ( .A(n745), .Q(n861) );
  BUF15 U490 ( .A(n112), .Q(n829) );
  OAI212 U491 ( .A(n5), .B(n46), .C(n47), .Q(n45) );
  AOI211 U493 ( .A(n877), .B(n190), .C(n191), .Q(n189) );
  NAND21 U494 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U495 ( .A(n151), .Q(n851) );
  XNR22 U498 ( .A(n7), .B(n41), .Q(SUM[31]) );
  OAI212 U503 ( .A(n42), .B(n830), .C(n43), .Q(n41) );
  NOR24 U504 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR21 U505 ( .A(n126), .B(n856), .Q(n122) );
  INV3 U506 ( .A(n53), .Q(n824) );
  NAND22 U507 ( .A(n111), .B(n55), .Q(n53) );
  INV3 U508 ( .A(n830), .Q(n825) );
  INV2 U509 ( .A(n830), .Q(n831) );
  NAND24 U511 ( .A(n592), .B(n65), .Q(n63) );
  NAND21 U512 ( .A(B[15]), .B(A[15]), .Q(n186) );
  NAND22 U513 ( .A(B[14]), .B(A[14]), .Q(n195) );
  NAND21 U514 ( .A(n111), .B(n853), .Q(n91) );
  AOI211 U515 ( .A(n829), .B(n853), .C(n98), .Q(n92) );
  NAND22 U517 ( .A(B[21]), .B(A[21]), .Q(n138) );
  NOR24 U518 ( .A(B[25]), .B(A[25]), .Q(n99) );
  OAI212 U520 ( .A(n830), .B(n82), .C(n83), .Q(n81) );
  NAND21 U521 ( .A(n111), .B(n840), .Q(n73) );
  XNR22 U522 ( .A(n9), .B(n63), .Q(SUM[29]) );
  AOI212 U523 ( .A(n183), .B(n204), .C(n184), .Q(n182) );
  NAND28 U524 ( .A(n77), .B(n853), .Q(n6) );
  NOR24 U525 ( .A(n79), .B(n88), .Q(n77) );
  XNR22 U527 ( .A(n11), .B(n81), .Q(SUM[27]) );
  OAI212 U528 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND24 U529 ( .A(n135), .B(n115), .Q(n113) );
  OAI212 U530 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  NOR23 U531 ( .A(n61), .B(n70), .Q(n59) );
  INV4 U532 ( .A(n70), .Q(n869) );
  CLKIN6 U533 ( .A(n59), .Q(n865) );
  NOR24 U534 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND21 U535 ( .A(n111), .B(n868), .Q(n102) );
  OAI211 U536 ( .A(n140), .B(n830), .C(n141), .Q(n139) );
  NOR23 U537 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND21 U538 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NOR24 U539 ( .A(B[22]), .B(A[22]), .Q(n126) );
  OAI212 U540 ( .A(n205), .B(n213), .C(n206), .Q(n204) );
  OAI211 U541 ( .A(n151), .B(n830), .C(n508), .Q(n146) );
  NAND22 U542 ( .A(B[23]), .B(A[23]), .Q(n118) );
  NAND24 U543 ( .A(n54), .B(n826), .Q(n52) );
  XNR22 U544 ( .A(n8), .B(n52), .Q(SUM[30]) );
  XOR20 U545 ( .A(n30), .B(n887), .Q(SUM[8]) );
  AOI212 U547 ( .A(n172), .B(n153), .C(n154), .Q(n508) );
  NAND20 U548 ( .A(n879), .B(n203), .Q(n197) );
  CLKIN0 U550 ( .A(n240), .Q(n884) );
  INV2 U551 ( .A(n255), .Q(n888) );
  INV1 U552 ( .A(n428), .Q(n847) );
  INV0 U553 ( .A(n239), .Q(n883) );
  AOI210 U554 ( .A(n877), .B(n203), .C(n204), .Q(n198) );
  CLKIN0 U555 ( .A(n163), .Q(n858) );
  INV0 U556 ( .A(n145), .Q(n863) );
  INV0 U557 ( .A(n231), .Q(n881) );
  INV0 U558 ( .A(n213), .Q(n876) );
  INV0 U559 ( .A(n244), .Q(n885) );
  INV0 U560 ( .A(n176), .Q(n849) );
  INV0 U561 ( .A(n241), .Q(n882) );
  INV0 U562 ( .A(n817), .Q(n873) );
  NOR22 U563 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR20 U564 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND21 U565 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND21 U566 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U567 ( .A(n39), .Q(n870) );
  NAND20 U568 ( .A(n888), .B(n256), .Q(n32) );
  INV3 U569 ( .A(n219), .Q(n879) );
  INV3 U570 ( .A(n171), .Q(n850) );
  AOI211 U571 ( .A(n829), .B(n837), .C(n85), .Q(n83) );
  INV3 U572 ( .A(n203), .Q(n874) );
  AOI211 U573 ( .A(n893), .B(n258), .C(n259), .Q(n257) );
  INV3 U574 ( .A(n268), .Q(n893) );
  NAND22 U575 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U576 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U577 ( .A(n252), .B(n255), .Q(n250) );
  AOI210 U578 ( .A(n848), .B(n862), .C(n863), .Q(n141) );
  NAND20 U579 ( .A(n171), .B(n859), .Q(n158) );
  AOI211 U580 ( .A(n428), .B(n859), .C(n858), .Q(n159) );
  AOI211 U581 ( .A(n829), .B(n868), .C(n867), .Q(n103) );
  NAND20 U582 ( .A(n239), .B(n880), .Q(n226) );
  AOI210 U583 ( .A(n240), .B(n880), .C(n881), .Q(n227) );
  NAND22 U584 ( .A(n879), .B(n190), .Q(n188) );
  NAND22 U585 ( .A(n879), .B(n875), .Q(n208) );
  INV3 U586 ( .A(n51), .Q(n834) );
  INV3 U587 ( .A(n230), .Q(n880) );
  INV3 U588 ( .A(n162), .Q(n859) );
  INV3 U589 ( .A(n212), .Q(n875) );
  NAND22 U590 ( .A(n886), .B(n253), .Q(n31) );
  INV3 U591 ( .A(n252), .Q(n886) );
  NAND22 U592 ( .A(n844), .B(n426), .Q(n580) );
  INV3 U593 ( .A(n61), .Q(n864) );
  INV3 U594 ( .A(n223), .Q(n878) );
  INV3 U595 ( .A(n265), .Q(n890) );
  NAND22 U596 ( .A(n892), .B(n272), .Q(n35) );
  INV3 U597 ( .A(n271), .Q(n892) );
  NAND22 U598 ( .A(n889), .B(n261), .Q(n33) );
  INV3 U599 ( .A(n260), .Q(n889) );
  INV3 U600 ( .A(n274), .Q(n894) );
  INV3 U601 ( .A(n278), .Q(n895) );
  AOI211 U602 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U603 ( .A(n271), .B(n274), .Q(n269) );
  NOR21 U604 ( .A(n260), .B(n265), .Q(n258) );
  INV3 U605 ( .A(n277), .Q(n896) );
  INV3 U606 ( .A(n266), .Q(n891) );
  NOR22 U607 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NAND22 U608 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND22 U609 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND22 U610 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND22 U611 ( .A(B[25]), .B(A[25]), .Q(n100) );
  NAND22 U612 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND22 U613 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NOR21 U614 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U615 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR21 U616 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U617 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR21 U618 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U619 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U620 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U621 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND22 U622 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND22 U623 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NOR21 U624 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U625 ( .A(n280), .Q(n898) );
  NOR21 U626 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U627 ( .A(A[0]), .B(B[0]), .Q(n281) );
  XNR21 U628 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND22 U629 ( .A(n870), .B(n40), .Q(n7) );
  NAND20 U630 ( .A(n100), .B(n854), .Q(n13) );
  NAND20 U631 ( .A(n838), .B(n89), .Q(n12) );
  NAND20 U632 ( .A(n864), .B(n62), .Q(n9) );
  XOR20 U633 ( .A(n22), .B(n830), .Q(SUM[16]) );
  NAND20 U634 ( .A(n849), .B(n177), .Q(n22) );
  XNR21 U635 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U636 ( .A(n880), .B(n231), .Q(n28) );
  XNR21 U637 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U638 ( .A(n878), .B(n224), .Q(n27) );
  XNR21 U639 ( .A(n24), .B(n196), .Q(SUM[14]) );
  NAND20 U640 ( .A(n195), .B(n871), .Q(n24) );
  XNR21 U641 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U642 ( .A(n873), .B(n206), .Q(n25) );
  NAND20 U643 ( .A(n885), .B(n245), .Q(n30) );
  XNR21 U644 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U645 ( .A(n882), .B(n242), .Q(n29) );
  XNR21 U646 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U647 ( .A(n832), .B(n186), .Q(n23) );
  XNR21 U648 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U649 ( .A(n875), .B(n213), .Q(n26) );
  NAND20 U650 ( .A(n860), .B(n174), .Q(n21) );
  XNR21 U651 ( .A(n17), .B(n139), .Q(SUM[21]) );
  NAND20 U652 ( .A(n138), .B(n855), .Q(n17) );
  XNR21 U653 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U654 ( .A(n857), .B(n156), .Q(n19) );
  XNR21 U655 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND20 U656 ( .A(n823), .B(n844), .Q(n16) );
  XNR21 U657 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND20 U658 ( .A(n861), .B(n118), .Q(n15) );
  XNR21 U659 ( .A(n18), .B(n146), .Q(SUM[20]) );
  NAND20 U660 ( .A(n862), .B(n145), .Q(n18) );
  XNR21 U661 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND20 U662 ( .A(n859), .B(n163), .Q(n20) );
  XNR21 U663 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND20 U664 ( .A(n868), .B(n107), .Q(n14) );
  XOR21 U665 ( .A(n36), .B(n896), .Q(SUM[2]) );
  NAND22 U666 ( .A(n894), .B(n275), .Q(n36) );
  XNR21 U667 ( .A(n34), .B(n893), .Q(SUM[4]) );
  NAND22 U668 ( .A(n890), .B(n266), .Q(n34) );
  XOR21 U669 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U670 ( .A(n893), .B(n890), .C(n891), .Q(n262) );
  XOR21 U671 ( .A(n32), .B(n257), .Q(SUM[6]) );
  XOR21 U672 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U673 ( .A(n895), .B(n279), .Q(n37) );
  XNR21 U674 ( .A(n35), .B(n273), .Q(SUM[3]) );
  INV3 U675 ( .A(n38), .Q(SUM[0]) );
  NAND22 U676 ( .A(n898), .B(n281), .Q(n38) );
  INV3 U677 ( .A(n111), .Q(n845) );
endmodule


module adder_8 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_8_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module reg_2 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31,
         n34, n49, n51, n53, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n55, n56, n57, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n52, n54, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392;

  DF3 Dout_reg_29_ ( .D(n60), .C(Clk), .Q(Dout[29]), .QN(n49) );
  DF3 Dout_reg_28_ ( .D(n61), .C(Clk), .Q(Dout[28]), .QN(n34) );
  DF3 Dout_reg_27_ ( .D(n62), .C(Clk), .Q(Dout[27]), .QN(n31) );
  DF3 Dout_reg_26_ ( .D(n63), .C(Clk), .Q(Dout[26]), .QN(n29) );
  DF3 Dout_reg_25_ ( .D(n64), .C(Clk), .Q(Dout[25]), .QN(n27) );
  DF3 Dout_reg_24_ ( .D(n65), .C(Clk), .Q(Dout[24]), .QN(n25) );
  DF3 Dout_reg_23_ ( .D(n66), .C(Clk), .Q(Dout[23]), .QN(n23) );
  DF3 Dout_reg_22_ ( .D(n67), .C(Clk), .Q(Dout[22]), .QN(n21) );
  DF3 Dout_reg_21_ ( .D(n68), .C(Clk), .Q(Dout[21]), .QN(n19) );
  DF3 Dout_reg_20_ ( .D(n69), .C(Clk), .Q(Dout[20]), .QN(n17) );
  DF3 Dout_reg_19_ ( .D(n70), .C(Clk), .Q(Dout[19]), .QN(n15) );
  DF3 Dout_reg_18_ ( .D(n71), .C(Clk), .Q(Dout[18]), .QN(n13) );
  DF3 Dout_reg_17_ ( .D(n72), .C(Clk), .Q(Dout[17]), .QN(n11) );
  DF3 Dout_reg_16_ ( .D(n73), .C(Clk), .Q(Dout[16]), .QN(n9) );
  DF3 Dout_reg_15_ ( .D(n74), .C(Clk), .Q(Dout[15]), .QN(n7) );
  DF3 Dout_reg_14_ ( .D(n75), .C(Clk), .Q(Dout[14]), .QN(n5) );
  DF3 Dout_reg_13_ ( .D(n87), .C(Clk), .Q(Dout[13]), .QN(n82) );
  DF3 Dout_reg_12_ ( .D(n88), .C(Clk), .Q(Dout[12]), .QN(n81) );
  DF3 Dout_reg_11_ ( .D(n89), .C(Clk), .Q(Dout[11]), .QN(n80) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n79) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n78) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n77) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n76) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n57) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n56) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n55) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n85) );
  DF3 Dout_reg_30_ ( .D(n59), .C(Clk), .Q(Dout[30]), .QN(n51) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n83) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n86) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n84) );
  DF3 Dout_reg_31_ ( .D(n58), .C(Clk), .Q(Dout[31]), .QN(n53) );
  OAI222 U3 ( .A(n84), .B(n357), .C(n359), .D(n362), .Q(n99) );
  OAI222 U4 ( .A(n85), .B(n357), .C(n358), .D(n363), .Q(n98) );
  OAI222 U5 ( .A(n86), .B(n357), .C(n52), .D(n364), .Q(n97) );
  OAI222 U6 ( .A(n55), .B(n357), .C(n359), .D(n365), .Q(n96) );
  OAI222 U7 ( .A(n56), .B(n357), .C(n358), .D(n366), .Q(n95) );
  OAI222 U8 ( .A(n57), .B(n357), .C(n52), .D(n368), .Q(n94) );
  OAI222 U9 ( .A(n76), .B(n357), .C(n359), .D(n367), .Q(n93) );
  OAI222 U10 ( .A(n77), .B(n357), .C(n358), .D(n374), .Q(n92) );
  OAI222 U11 ( .A(n78), .B(n357), .C(n52), .D(n375), .Q(n91) );
  OAI222 U12 ( .A(n79), .B(n357), .C(n359), .D(n369), .Q(n90) );
  OAI222 U13 ( .A(n80), .B(n357), .C(n358), .D(n370), .Q(n89) );
  OAI222 U14 ( .A(n81), .B(n357), .C(n52), .D(n376), .Q(n88) );
  OAI222 U15 ( .A(n82), .B(n357), .C(n359), .D(n371), .Q(n87) );
  OAI222 U16 ( .A(n5), .B(n357), .C(n358), .D(n372), .Q(n75) );
  OAI222 U17 ( .A(n7), .B(n357), .C(n52), .D(n373), .Q(n74) );
  OAI222 U18 ( .A(n9), .B(n357), .C(n359), .D(n378), .Q(n73) );
  OAI222 U19 ( .A(n11), .B(n357), .C(n358), .D(n377), .Q(n72) );
  OAI222 U20 ( .A(n13), .B(n357), .C(n52), .D(n391), .Q(n71) );
  OAI222 U21 ( .A(n15), .B(n357), .C(n359), .D(n390), .Q(n70) );
  OAI222 U22 ( .A(n17), .B(n357), .C(n358), .D(n389), .Q(n69) );
  OAI222 U23 ( .A(n19), .B(n357), .C(n52), .D(n388), .Q(n68) );
  OAI222 U24 ( .A(n21), .B(n357), .C(n359), .D(n387), .Q(n67) );
  OAI222 U25 ( .A(n23), .B(n357), .C(n358), .D(n392), .Q(n66) );
  OAI222 U26 ( .A(n25), .B(n357), .C(n52), .D(n386), .Q(n65) );
  OAI222 U27 ( .A(n27), .B(n357), .C(n359), .D(n385), .Q(n64) );
  OAI222 U28 ( .A(n29), .B(n357), .C(n358), .D(n384), .Q(n63) );
  OAI222 U29 ( .A(n31), .B(n357), .C(n52), .D(n383), .Q(n62) );
  OAI222 U30 ( .A(n34), .B(n357), .C(n359), .D(n382), .Q(n61) );
  OAI222 U31 ( .A(n49), .B(n357), .C(n358), .D(n381), .Q(n60) );
  OAI222 U32 ( .A(n51), .B(n357), .C(n52), .D(n380), .Q(n59) );
  OAI222 U33 ( .A(n53), .B(n357), .C(n359), .D(n379), .Q(n58) );
  OAI222 U34 ( .A(n83), .B(n357), .C(n358), .D(n361), .Q(n100) );
  CLKIN3 U35 ( .A(Din[16]), .Q(n378) );
  CLKIN3 U36 ( .A(Din[31]), .Q(n379) );
  CLKIN3 U37 ( .A(Din[17]), .Q(n377) );
  CLKIN3 U38 ( .A(Din[19]), .Q(n390) );
  CLKIN3 U39 ( .A(Din[20]), .Q(n389) );
  CLKIN3 U40 ( .A(Din[22]), .Q(n387) );
  CLKIN3 U41 ( .A(Din[23]), .Q(n392) );
  CLKIN3 U42 ( .A(Din[25]), .Q(n385) );
  CLKIN3 U43 ( .A(Din[26]), .Q(n384) );
  CLKIN3 U44 ( .A(Din[28]), .Q(n382) );
  CLKIN3 U45 ( .A(Din[29]), .Q(n381) );
  CLKIN3 U46 ( .A(Din[30]), .Q(n380) );
  CLKIN3 U47 ( .A(Din[18]), .Q(n391) );
  CLKIN3 U48 ( .A(Din[21]), .Q(n388) );
  CLKIN3 U49 ( .A(Din[24]), .Q(n386) );
  CLKIN3 U50 ( .A(Din[27]), .Q(n383) );
  NAND22 U51 ( .A(n360), .B(n357), .Q(n359) );
  NAND22 U52 ( .A(n360), .B(n357), .Q(n358) );
  NAND22 U53 ( .A(n360), .B(n357), .Q(n52) );
  INV3 U54 ( .A(Reset), .Q(n360) );
  INV3 U55 ( .A(n54), .Q(n357) );
  INV3 U56 ( .A(Din[8]), .Q(n374) );
  INV3 U57 ( .A(Din[6]), .Q(n368) );
  INV3 U58 ( .A(Din[5]), .Q(n366) );
  INV3 U59 ( .A(Din[7]), .Q(n367) );
  INV3 U60 ( .A(Din[9]), .Q(n375) );
  INV3 U61 ( .A(Din[10]), .Q(n369) );
  INV3 U62 ( .A(Din[11]), .Q(n370) );
  INV3 U63 ( .A(Din[12]), .Q(n376) );
  INV3 U64 ( .A(Din[13]), .Q(n371) );
  INV3 U65 ( .A(Din[14]), .Q(n372) );
  INV3 U66 ( .A(Din[15]), .Q(n373) );
  INV3 U67 ( .A(Din[4]), .Q(n365) );
  INV3 U68 ( .A(Din[2]), .Q(n363) );
  INV3 U69 ( .A(Din[0]), .Q(n361) );
  INV3 U70 ( .A(Din[3]), .Q(n364) );
  INV3 U71 ( .A(Din[1]), .Q(n362) );
  NOR21 U72 ( .A(Load), .B(Reset), .Q(n54) );
endmodule


module reg_1 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n3, n5, n7, n9, n11, n13, n17, n19, n21, n23, n25, n27, n29, n31, n34,
         n49, n51, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n68,
         n69, n70, n71, n72, n73, n55, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394;

  DF3 Dout_reg_15_ ( .D(n72), .C(Clk), .Q(Dout[15]), .QN(n5) );
  DF3 Dout_reg_14_ ( .D(n73), .C(Clk), .Q(Dout[14]), .QN(n3) );
  DF3 Dout_reg_13_ ( .D(n87), .C(Clk), .Q(Dout[13]), .QN(n77) );
  DF3 Dout_reg_12_ ( .D(n88), .C(Clk), .Q(Dout[12]), .QN(n78) );
  DF3 Dout_reg_11_ ( .D(n89), .C(Clk), .Q(Dout[11]), .QN(n76) );
  DF3 Dout_reg_10_ ( .D(n90), .C(Clk), .Q(Dout[10]), .QN(n75) );
  DF3 Dout_reg_7_ ( .D(n93), .C(Clk), .Q(Dout[7]), .QN(n82) );
  DF3 Dout_reg_6_ ( .D(n94), .C(Clk), .Q(Dout[6]), .QN(n79) );
  DF3 Dout_reg_4_ ( .D(n96), .C(Clk), .Q(Dout[4]), .QN(n81) );
  DF3 Dout_reg_3_ ( .D(n97), .C(Clk), .Q(Dout[3]), .QN(n85) );
  DF3 Dout_reg_2_ ( .D(n98), .C(Clk), .Q(Dout[2]), .QN(n83) );
  DF3 Dout_reg_0_ ( .D(n100), .C(Clk), .Q(Dout[0]), .QN(n86) );
  DF3 Dout_reg_5_ ( .D(n95), .C(Clk), .Q(Dout[5]), .QN(n80) );
  DF3 Dout_reg_16_ ( .D(n71), .C(Clk), .Q(Dout[16]), .QN(n7) );
  DF3 Dout_reg_1_ ( .D(n99), .C(Clk), .Q(Dout[1]), .QN(n84) );
  DF3 Dout_reg_17_ ( .D(n70), .C(Clk), .Q(Dout[17]), .QN(n9) );
  DF3 Dout_reg_8_ ( .D(n92), .C(Clk), .Q(Dout[8]), .QN(n55) );
  DF3 Dout_reg_18_ ( .D(n69), .C(Clk), .Q(Dout[18]), .QN(n11) );
  DF3 Dout_reg_24_ ( .D(n63), .C(Clk), .Q(Dout[24]), .QN(n23) );
  DF3 Dout_reg_23_ ( .D(n64), .C(Clk), .Q(Dout[23]), .QN(n21) );
  DF3 Dout_reg_21_ ( .D(n66), .C(Clk), .Q(Dout[21]), .QN(n17) );
  DF3 Dout_reg_19_ ( .D(n68), .C(Clk), .Q(Dout[19]), .QN(n13) );
  OAI222 U3 ( .A(n103), .B(n359), .C(n361), .D(n394), .Q(n104) );
  OAI222 U4 ( .A(n84), .B(n359), .C(n360), .D(n364), .Q(n99) );
  OAI222 U5 ( .A(n83), .B(n359), .C(n101), .D(n366), .Q(n98) );
  OAI222 U6 ( .A(n85), .B(n359), .C(n361), .D(n365), .Q(n97) );
  OAI222 U7 ( .A(n81), .B(n359), .C(n360), .D(n367), .Q(n96) );
  OAI222 U8 ( .A(n80), .B(n359), .C(n101), .D(n368), .Q(n95) );
  OAI222 U9 ( .A(n79), .B(n359), .C(n361), .D(n370), .Q(n94) );
  OAI222 U10 ( .A(n82), .B(n359), .C(n360), .D(n369), .Q(n93) );
  OAI222 U11 ( .A(n55), .B(n359), .C(n101), .D(n378), .Q(n92) );
  OAI222 U12 ( .A(n74), .B(n359), .C(n361), .D(n377), .Q(n91) );
  OAI222 U13 ( .A(n75), .B(n359), .C(n360), .D(n375), .Q(n90) );
  OAI222 U14 ( .A(n76), .B(n359), .C(n101), .D(n374), .Q(n89) );
  OAI222 U15 ( .A(n78), .B(n359), .C(n376), .D(n361), .Q(n88) );
  OAI222 U16 ( .A(n77), .B(n359), .C(n360), .D(n371), .Q(n87) );
  OAI222 U17 ( .A(n3), .B(n359), .C(n101), .D(n373), .Q(n73) );
  OAI222 U18 ( .A(n5), .B(n359), .C(n361), .D(n372), .Q(n72) );
  OAI222 U19 ( .A(n7), .B(n359), .C(n360), .D(n383), .Q(n71) );
  OAI222 U20 ( .A(n9), .B(n359), .C(n101), .D(n392), .Q(n70) );
  OAI222 U21 ( .A(n11), .B(n359), .C(n361), .D(n390), .Q(n69) );
  OAI222 U22 ( .A(n13), .B(n359), .C(n360), .D(n386), .Q(n68) );
  OAI222 U23 ( .A(n17), .B(n359), .C(n101), .D(n391), .Q(n66) );
  OAI222 U24 ( .A(n19), .B(n359), .C(n361), .D(n393), .Q(n65) );
  OAI222 U25 ( .A(n21), .B(n359), .C(n360), .D(n384), .Q(n64) );
  OAI222 U26 ( .A(n23), .B(n359), .C(n101), .D(n385), .Q(n63) );
  OAI222 U27 ( .A(n25), .B(n359), .C(n361), .D(n388), .Q(n62) );
  OAI222 U28 ( .A(n27), .B(n359), .C(n360), .D(n382), .Q(n61) );
  OAI222 U29 ( .A(n29), .B(n359), .C(n381), .D(n101), .Q(n60) );
  OAI222 U30 ( .A(n31), .B(n359), .C(n361), .D(n389), .Q(n59) );
  OAI222 U31 ( .A(n34), .B(n359), .C(n360), .D(n380), .Q(n58) );
  OAI222 U32 ( .A(n49), .B(n359), .C(n379), .D(n101), .Q(n57) );
  OAI222 U33 ( .A(n51), .B(n359), .C(n361), .D(n387), .Q(n56) );
  OAI222 U34 ( .A(n86), .B(n359), .C(n360), .D(n363), .Q(n100) );
  DF1 Dout_reg_22_ ( .D(n65), .C(Clk), .Q(Dout[22]), .QN(n19) );
  DF1 Dout_reg_30_ ( .D(n57), .C(Clk), .Q(Dout[30]), .QN(n49) );
  DF1 Dout_reg_27_ ( .D(n60), .C(Clk), .Q(Dout[27]), .QN(n29) );
  DF1 Dout_reg_31_ ( .D(n56), .C(Clk), .Q(Dout[31]), .QN(n51) );
  DF1 Dout_reg_29_ ( .D(n58), .C(Clk), .Q(Dout[29]), .QN(n34) );
  DF1 Dout_reg_20_ ( .D(n104), .C(Clk), .Q(Dout[20]), .QN(n103) );
  DF3 Dout_reg_9_ ( .D(n91), .C(Clk), .Q(Dout[9]), .QN(n74) );
  DF3 Dout_reg_26_ ( .D(n61), .C(Clk), .Q(Dout[26]), .QN(n27) );
  DF3 Dout_reg_28_ ( .D(n59), .C(Clk), .Q(Dout[28]), .QN(n31) );
  DF3 Dout_reg_25_ ( .D(n62), .C(Clk), .Q(Dout[25]), .QN(n25) );
  INV3 U35 ( .A(Din[25]), .Q(n388) );
  INV3 U36 ( .A(Din[28]), .Q(n389) );
  INV3 U37 ( .A(Din[20]), .Q(n394) );
  INV3 U38 ( .A(Din[27]), .Q(n381) );
  INV3 U39 ( .A(Din[31]), .Q(n387) );
  INV3 U40 ( .A(Din[29]), .Q(n380) );
  INV3 U41 ( .A(Din[30]), .Q(n379) );
  INV3 U42 ( .A(Din[23]), .Q(n384) );
  INV3 U43 ( .A(Din[26]), .Q(n382) );
  INV3 U44 ( .A(Din[12]), .Q(n376) );
  INV3 U45 ( .A(Din[17]), .Q(n392) );
  INV3 U46 ( .A(Din[9]), .Q(n377) );
  CLKIN3 U47 ( .A(Din[8]), .Q(n378) );
  INV2 U48 ( .A(Din[22]), .Q(n393) );
  INV2 U49 ( .A(Din[19]), .Q(n386) );
  INV2 U50 ( .A(Din[18]), .Q(n390) );
  INV2 U51 ( .A(Din[16]), .Q(n383) );
  INV2 U52 ( .A(Din[13]), .Q(n371) );
  INV2 U53 ( .A(Din[15]), .Q(n372) );
  INV2 U54 ( .A(Din[10]), .Q(n375) );
  INV2 U55 ( .A(Din[24]), .Q(n385) );
  INV2 U56 ( .A(Din[21]), .Q(n391) );
  INV2 U57 ( .A(Din[14]), .Q(n373) );
  INV2 U58 ( .A(Din[11]), .Q(n374) );
  CLKIN3 U59 ( .A(Din[7]), .Q(n369) );
  NAND22 U60 ( .A(n362), .B(n359), .Q(n360) );
  NAND22 U61 ( .A(n362), .B(n359), .Q(n361) );
  NAND22 U62 ( .A(n362), .B(n359), .Q(n101) );
  INV3 U63 ( .A(Reset), .Q(n362) );
  INV3 U64 ( .A(n102), .Q(n359) );
  INV3 U65 ( .A(Din[3]), .Q(n365) );
  INV3 U66 ( .A(Din[5]), .Q(n368) );
  INV3 U67 ( .A(Din[6]), .Q(n370) );
  INV3 U68 ( .A(Din[1]), .Q(n364) );
  INV3 U69 ( .A(Din[4]), .Q(n367) );
  INV3 U70 ( .A(Din[2]), .Q(n366) );
  INV3 U71 ( .A(Din[0]), .Q(n363) );
  NOR21 U72 ( .A(Load), .B(Reset), .Q(n102) );
endmodule


module adder_7_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n212, n213, n214, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n232, n239, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n422, n423,
         n556, n557, n694, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827;

  OAI212 U43 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U101 ( .A(n794), .B(n762), .C(n797), .Q(n108) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n762), .C(n121), .Q(n119) );
  OAI212 U141 ( .A(n140), .B(n762), .C(n141), .Q(n139) );
  OAI212 U165 ( .A(n158), .B(n762), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n792), .B(n762), .C(n795), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U189 ( .A(n176), .B(n762), .C(n177), .Q(n175) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  AOI212 U321 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  AOI212 U349 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  OAI212 U353 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U379 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U421 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U618 ( .A(n274), .B(n785), .C(n275), .Q(n273) );
  OAI212 U431 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  OAI212 U474 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  AOI212 U487 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U373 ( .A(n789), .B(n776), .C(n790), .Q(n232) );
  OAI212 U381 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  OAI212 U424 ( .A(n194), .B(n768), .C(n195), .Q(n191) );
  OAI212 U433 ( .A(n64), .B(n762), .C(n65), .Q(n63) );
  OAI212 U472 ( .A(n88), .B(n805), .C(n89), .Q(n85) );
  OAI212 U375 ( .A(n268), .B(n248), .C(n249), .Q(n556) );
  OAI212 U417 ( .A(n244), .B(n776), .C(n245), .Q(n243) );
  OAI212 U456 ( .A(n188), .B(n776), .C(n189), .Q(n187) );
  OAI212 U515 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U382 ( .A(n226), .B(n776), .C(n227), .Q(n225) );
  AOI212 U442 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U380 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U392 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U412 ( .A(n208), .B(n776), .C(n209), .Q(n207) );
  OAI212 U419 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U355 ( .A(n275), .B(n271), .C(n272), .Q(n694) );
  OAI212 U404 ( .A(n268), .B(n248), .C(n249), .Q(n247) );
  OAI212 U405 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI212 U426 ( .A(n53), .B(n762), .C(n54), .Q(n52) );
  OAI212 U437 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U448 ( .A(n129), .B(n762), .C(n130), .Q(n128) );
  OAI212 U458 ( .A(n82), .B(n762), .C(n83), .Q(n81) );
  AOI212 U464 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  XNR22 U350 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NOR23 U351 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NAND22 U352 ( .A(n239), .B(n221), .Q(n219) );
  INV2 U354 ( .A(n220), .Q(n773) );
  XNR22 U356 ( .A(n18), .B(n146), .Q(SUM[20]) );
  XOR22 U357 ( .A(n22), .B(n762), .Q(SUM[16]) );
  NOR22 U358 ( .A(n260), .B(n265), .Q(n258) );
  NOR22 U359 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NOR23 U360 ( .A(n117), .B(n126), .Q(n115) );
  NOR22 U361 ( .A(B[23]), .B(A[23]), .Q(n117) );
  XNR22 U362 ( .A(n24), .B(n196), .Q(SUM[14]) );
  XNR22 U363 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NOR21 U364 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR22 U365 ( .A(n252), .B(n255), .Q(n250) );
  NOR22 U366 ( .A(B[22]), .B(A[22]), .Q(n126) );
  INV3 U367 ( .A(n152), .Q(n796) );
  NOR22 U368 ( .A(n271), .B(n274), .Q(n269) );
  NOR22 U369 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR22 U370 ( .A(n223), .B(n230), .Q(n221) );
  NAND24 U371 ( .A(n203), .B(n183), .Q(n181) );
  NAND23 U372 ( .A(n258), .B(n250), .Q(n248) );
  NOR21 U374 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR23 U376 ( .A(B[1]), .B(A[1]), .Q(n278) );
  XNR21 U377 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI212 U378 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI211 U383 ( .A(n197), .B(n776), .C(n198), .Q(n196) );
  NAND22 U384 ( .A(n793), .B(n822), .Q(n140) );
  INV3 U385 ( .A(n144), .Q(n822) );
  OAI210 U386 ( .A(n42), .B(n762), .C(n43), .Q(n41) );
  NAND22 U387 ( .A(n59), .B(n823), .Q(n46) );
  XNR22 U388 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND22 U389 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND21 U390 ( .A(n822), .B(n145), .Q(n18) );
  OAI210 U391 ( .A(n126), .B(n812), .C(n127), .Q(n123) );
  INV1 U393 ( .A(n277), .Q(n785) );
  XNR22 U394 ( .A(n26), .B(n214), .Q(SUM[12]) );
  AOI212 U395 ( .A(n112), .B(n84), .C(n85), .Q(n83) );
  AOI212 U396 ( .A(n112), .B(n97), .C(n98), .Q(n92) );
  AOI211 U397 ( .A(n112), .B(n809), .C(n806), .Q(n74) );
  NOR24 U398 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NAND21 U399 ( .A(A[25]), .B(B[25]), .Q(n100) );
  OAI211 U400 ( .A(n73), .B(n762), .C(n74), .Q(n72) );
  NOR22 U401 ( .A(n79), .B(n88), .Q(n77) );
  NAND22 U402 ( .A(n111), .B(n66), .Q(n64) );
  NOR20 U403 ( .A(n70), .B(n6), .Q(n66) );
  NOR21 U406 ( .A(n126), .B(n814), .Q(n122) );
  NAND24 U407 ( .A(n135), .B(n115), .Q(n113) );
  XNR22 U408 ( .A(n13), .B(n101), .Q(SUM[25]) );
  XNR22 U409 ( .A(n14), .B(n108), .Q(SUM[24]) );
  NAND21 U410 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NOR24 U411 ( .A(n181), .B(n219), .Q(n179) );
  NOR22 U413 ( .A(n185), .B(n194), .Q(n183) );
  INV8 U414 ( .A(n556), .Q(n776) );
  NOR24 U415 ( .A(B[3]), .B(A[3]), .Q(n271) );
  XNR22 U416 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND22 U418 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND21 U420 ( .A(A[11]), .B(B[11]), .Q(n224) );
  BUF15 U422 ( .A(n178), .Q(n762) );
  AOI211 U423 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND22 U425 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NOR22 U427 ( .A(n241), .B(n244), .Q(n239) );
  NOR24 U428 ( .A(n113), .B(n151), .Q(n111) );
  NOR22 U429 ( .A(n155), .B(n162), .Q(n153) );
  INV0 U430 ( .A(n252), .Q(n777) );
  XNR22 U432 ( .A(n29), .B(n243), .Q(SUM[9]) );
  OAI211 U434 ( .A(n91), .B(n762), .C(n92), .Q(n90) );
  NAND21 U435 ( .A(n111), .B(n97), .Q(n91) );
  NOR23 U436 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND24 U438 ( .A(n422), .B(n423), .Q(SUM[17]) );
  NOR23 U439 ( .A(n205), .B(n212), .Q(n203) );
  NOR22 U440 ( .A(B[12]), .B(A[12]), .Q(n212) );
  INV3 U441 ( .A(n203), .Q(n767) );
  AOI211 U443 ( .A(n269), .B(n277), .C(n694), .Q(n557) );
  XNR22 U444 ( .A(n17), .B(n139), .Q(SUM[21]) );
  XNR22 U445 ( .A(n23), .B(n187), .Q(SUM[15]) );
  OAI211 U446 ( .A(n102), .B(n762), .C(n103), .Q(n101) );
  OAI212 U447 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  AOI212 U449 ( .A(n781), .B(n258), .C(n259), .Q(n257) );
  XNR22 U450 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U451 ( .A(n769), .B(n213), .Q(n26) );
  INV0 U452 ( .A(n213), .Q(n770) );
  XOR20 U453 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NOR23 U454 ( .A(B[10]), .B(A[10]), .Q(n230) );
  OAI211 U455 ( .A(n219), .B(n776), .C(n220), .Q(n214) );
  XNR22 U457 ( .A(n15), .B(n119), .Q(SUM[23]) );
  NAND21 U459 ( .A(A[17]), .B(B[17]), .Q(n174) );
  AOI211 U460 ( .A(n796), .B(n822), .C(n821), .Q(n141) );
  NAND21 U461 ( .A(n793), .B(n122), .Q(n120) );
  NAND22 U462 ( .A(n793), .B(n135), .Q(n129) );
  INV3 U463 ( .A(n151), .Q(n793) );
  CLKIN1 U465 ( .A(n97), .Q(n808) );
  INV1 U466 ( .A(n6), .Q(n809) );
  CLKIN0 U467 ( .A(n204), .Q(n768) );
  NAND21 U468 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND21 U469 ( .A(A[15]), .B(B[15]), .Q(n186) );
  AOI211 U470 ( .A(n773), .B(n190), .C(n191), .Q(n189) );
  INV2 U471 ( .A(n557), .Q(n781) );
  INV0 U473 ( .A(n231), .Q(n775) );
  INV2 U475 ( .A(n98), .Q(n805) );
  NAND20 U476 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND20 U477 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND21 U478 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U479 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND21 U480 ( .A(A[22]), .B(B[22]), .Q(n127) );
  CLKIN3 U481 ( .A(n60), .Q(n818) );
  AOI211 U482 ( .A(n773), .B(n203), .C(n204), .Q(n198) );
  NAND22 U483 ( .A(n772), .B(n203), .Q(n197) );
  CLKIN0 U484 ( .A(n240), .Q(n790) );
  NAND21 U485 ( .A(n771), .B(n224), .Q(n27) );
  NAND21 U486 ( .A(n788), .B(n242), .Q(n29) );
  CLKIN0 U488 ( .A(n112), .Q(n797) );
  INV0 U489 ( .A(n106), .Q(n807) );
  NAND20 U490 ( .A(n791), .B(n177), .Q(n22) );
  NAND20 U491 ( .A(n819), .B(n71), .Q(n10) );
  NAND20 U492 ( .A(n782), .B(n272), .Q(n35) );
  NAND21 U493 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND22 U494 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND22 U495 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NOR20 U496 ( .A(n820), .B(n6), .Q(n55) );
  NAND20 U497 ( .A(n111), .B(n807), .Q(n102) );
  NAND21 U498 ( .A(n111), .B(n84), .Q(n82) );
  OAI210 U499 ( .A(n820), .B(n5), .C(n818), .Q(n56) );
  INV1 U500 ( .A(n5), .Q(n806) );
  CLKIN0 U501 ( .A(n172), .Q(n795) );
  NOR20 U502 ( .A(n46), .B(n6), .Q(n44) );
  NAND21 U503 ( .A(n772), .B(n190), .Q(n188) );
  NAND20 U504 ( .A(n239), .B(n774), .Q(n226) );
  NAND20 U505 ( .A(n171), .B(n802), .Q(n158) );
  CLKIN3 U506 ( .A(n59), .Q(n820) );
  CLKIN0 U507 ( .A(n239), .Q(n789) );
  NOR22 U508 ( .A(n99), .B(n106), .Q(n97) );
  NOR22 U509 ( .A(n137), .B(n144), .Q(n135) );
  INV0 U510 ( .A(n176), .Q(n791) );
  CLKIN0 U511 ( .A(n126), .Q(n811) );
  CLKIN0 U512 ( .A(n171), .Q(n792) );
  NAND20 U513 ( .A(n802), .B(n163), .Q(n20) );
  INV0 U514 ( .A(n255), .Q(n778) );
  INV0 U516 ( .A(n99), .Q(n817) );
  INV0 U517 ( .A(n79), .Q(n826) );
  INV0 U518 ( .A(n70), .Q(n819) );
  INV0 U519 ( .A(n205), .Q(n766) );
  INV0 U520 ( .A(n155), .Q(n815) );
  INV0 U521 ( .A(n117), .Q(n810) );
  NAND20 U522 ( .A(n779), .B(n266), .Q(n34) );
  INV0 U523 ( .A(n223), .Q(n771) );
  AOI210 U524 ( .A(n60), .B(n823), .C(n824), .Q(n47) );
  INV0 U525 ( .A(n244), .Q(n801) );
  INV0 U526 ( .A(n260), .Q(n787) );
  INV0 U527 ( .A(n173), .Q(n800) );
  INV0 U528 ( .A(n241), .Q(n788) );
  NAND20 U529 ( .A(n774), .B(n231), .Q(n28) );
  INV0 U530 ( .A(n185), .Q(n763) );
  XOR20 U531 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND20 U532 ( .A(n798), .B(n279), .Q(n37) );
  NAND20 U533 ( .A(n783), .B(n275), .Q(n36) );
  INV0 U534 ( .A(n274), .Q(n783) );
  INV0 U535 ( .A(n271), .Q(n782) );
  INV0 U536 ( .A(n266), .Q(n780) );
  NOR22 U537 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NOR22 U538 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND20 U539 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND21 U540 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NAND21 U541 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND20 U542 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND21 U543 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NAND20 U544 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND21 U545 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND22 U546 ( .A(n111), .B(n809), .Q(n73) );
  INV3 U547 ( .A(n111), .Q(n794) );
  NAND20 U548 ( .A(n111), .B(n44), .Q(n42) );
  INV3 U549 ( .A(n219), .Q(n772) );
  NAND22 U550 ( .A(n97), .B(n77), .Q(n6) );
  NAND22 U551 ( .A(n171), .B(n153), .Q(n151) );
  AOI210 U552 ( .A(n796), .B(n135), .C(n136), .Q(n130) );
  NAND22 U553 ( .A(n799), .B(n764), .Q(n423) );
  INV3 U554 ( .A(n21), .Q(n799) );
  NAND22 U555 ( .A(n772), .B(n769), .Q(n208) );
  NAND22 U556 ( .A(n810), .B(n118), .Q(n15) );
  XNR21 U557 ( .A(n11), .B(n81), .Q(SUM[27]) );
  NAND22 U558 ( .A(n826), .B(n80), .Q(n11) );
  NAND22 U559 ( .A(n813), .B(n138), .Q(n17) );
  INV3 U560 ( .A(n137), .Q(n813) );
  XOR21 U561 ( .A(n30), .B(n776), .Q(SUM[8]) );
  NAND22 U562 ( .A(n801), .B(n245), .Q(n30) );
  NAND22 U563 ( .A(n778), .B(n256), .Q(n32) );
  INV3 U564 ( .A(n51), .Q(n824) );
  XNR21 U565 ( .A(n254), .B(n31), .Q(SUM[7]) );
  NAND22 U566 ( .A(n777), .B(n253), .Q(n31) );
  NAND22 U567 ( .A(n816), .B(n89), .Q(n12) );
  INV3 U568 ( .A(n88), .Q(n816) );
  XNR21 U569 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR21 U570 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NAND22 U571 ( .A(n827), .B(n62), .Q(n9) );
  INV3 U572 ( .A(n61), .Q(n827) );
  NAND22 U573 ( .A(n807), .B(n107), .Q(n14) );
  XNR21 U574 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND22 U575 ( .A(n811), .B(n127), .Q(n16) );
  XNR21 U576 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NAND22 U577 ( .A(n823), .B(n51), .Q(n8) );
  NAND20 U578 ( .A(n111), .B(n55), .Q(n53) );
  NOR21 U579 ( .A(n173), .B(n176), .Q(n171) );
  NOR21 U580 ( .A(n61), .B(n70), .Q(n59) );
  INV3 U581 ( .A(n107), .Q(n804) );
  NAND22 U582 ( .A(n817), .B(n100), .Q(n13) );
  NAND22 U583 ( .A(n815), .B(n156), .Q(n19) );
  NAND22 U584 ( .A(n766), .B(n206), .Q(n25) );
  NAND22 U585 ( .A(n765), .B(n195), .Q(n24) );
  INV3 U586 ( .A(n194), .Q(n765) );
  NAND22 U587 ( .A(n763), .B(n186), .Q(n23) );
  NOR21 U588 ( .A(n88), .B(n808), .Q(n84) );
  INV0 U589 ( .A(n135), .Q(n814) );
  AOI210 U590 ( .A(n172), .B(n802), .C(n803), .Q(n159) );
  INV3 U591 ( .A(n163), .Q(n803) );
  AOI211 U592 ( .A(n796), .B(n122), .C(n123), .Q(n121) );
  INV0 U593 ( .A(n136), .Q(n812) );
  INV3 U594 ( .A(n145), .Q(n821) );
  AOI211 U595 ( .A(n773), .B(n769), .C(n770), .Q(n209) );
  NAND22 U596 ( .A(n800), .B(n174), .Q(n21) );
  INV3 U597 ( .A(n162), .Q(n802) );
  INV3 U598 ( .A(n212), .Q(n769) );
  INV3 U599 ( .A(n230), .Q(n774) );
  NOR21 U600 ( .A(n194), .B(n767), .Q(n190) );
  XOR21 U601 ( .A(n33), .B(n262), .Q(SUM[5]) );
  NAND22 U602 ( .A(n787), .B(n261), .Q(n33) );
  AOI210 U603 ( .A(n781), .B(n779), .C(n780), .Q(n262) );
  XOR21 U604 ( .A(n36), .B(n785), .Q(SUM[2]) );
  XNR21 U605 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XNR20 U606 ( .A(n34), .B(n781), .Q(SUM[4]) );
  INV3 U607 ( .A(n278), .Q(n798) );
  INV3 U608 ( .A(n265), .Q(n779) );
  NOR21 U609 ( .A(B[28]), .B(A[28]), .Q(n70) );
  XNR21 U610 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U611 ( .A(n825), .B(n40), .Q(n7) );
  NAND22 U612 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR22 U613 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR22 U614 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR22 U615 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR22 U616 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR22 U617 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR22 U619 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR22 U620 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR22 U621 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR22 U622 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR22 U623 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR22 U624 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR22 U625 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR21 U626 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND22 U627 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U628 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND22 U629 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U630 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND22 U631 ( .A(B[1]), .B(A[1]), .Q(n279) );
  INV3 U632 ( .A(n50), .Q(n823) );
  NOR21 U633 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NAND22 U634 ( .A(A[30]), .B(B[30]), .Q(n51) );
  INV3 U635 ( .A(n39), .Q(n825) );
  NOR21 U636 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U637 ( .A(n38), .Q(SUM[0]) );
  NAND20 U638 ( .A(n786), .B(n281), .Q(n38) );
  INV3 U639 ( .A(n280), .Q(n786) );
  NOR20 U640 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U641 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND22 U642 ( .A(n21), .B(n175), .Q(n422) );
  INV3 U643 ( .A(n175), .Q(n764) );
  AOI210 U644 ( .A(n112), .B(n44), .C(n45), .Q(n43) );
  AOI210 U645 ( .A(n112), .B(n55), .C(n56), .Q(n54) );
  AOI210 U646 ( .A(n112), .B(n66), .C(n67), .Q(n65) );
  AOI211 U647 ( .A(n112), .B(n807), .C(n804), .Q(n103) );
  OAI211 U648 ( .A(n151), .B(n762), .C(n152), .Q(n146) );
  AOI210 U649 ( .A(n240), .B(n774), .C(n775), .Q(n227) );
endmodule


module adder_7 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_7_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n48, n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n69, n70, n71, n72, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n99, n100,
         n101, n102, n103, n106, n107, n108, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n127, n128, n129, n130,
         n131, n132, n137, n138, n139, n140, n141, n144, n145, n146, n147,
         n148, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n167, n168, n173, n174, n175, n176, n177, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n195,
         n196, n197, n198, n199, n200, n205, n206, n207, n208, n209, n212,
         n213, n214, n215, n216, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n235, n236, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n737, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800;

  OAI212 U15 ( .A(n44), .B(n76), .C(n45), .Q(n43) );
  OAI212 U29 ( .A(n747), .B(n76), .C(n748), .Q(n54) );
  OAI212 U33 ( .A(n69), .B(n59), .C(n60), .Q(n58) );
  OAI212 U43 ( .A(n66), .B(n76), .C(n69), .Q(n65) );
  OAI212 U59 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U69 ( .A(n86), .B(n756), .C(n89), .Q(n85) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n94) );
  OAI212 U105 ( .A(n113), .B(n148), .C(n114), .Q(n3) );
  OAI212 U115 ( .A(n120), .B(n737), .C(n121), .Q(n119) );
  OAI212 U119 ( .A(n124), .B(n765), .C(n127), .Q(n123) );
  OAI212 U127 ( .A(n129), .B(n737), .C(n130), .Q(n128) );
  OAI212 U135 ( .A(n145), .B(n137), .C(n138), .Q(n132) );
  OAI212 U141 ( .A(n140), .B(n737), .C(n141), .Q(n139) );
  OAI212 U151 ( .A(n147), .B(n737), .C(n148), .Q(n146) );
  OAI212 U159 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U165 ( .A(n158), .B(n737), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n774), .B(n737), .C(n775), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n168) );
  OAI212 U197 ( .A(n181), .B(n216), .C(n182), .Q(n180) );
  OAI212 U201 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI212 U207 ( .A(n188), .B(n742), .C(n189), .Q(n187) );
  OAI212 U211 ( .A(n192), .B(n779), .C(n195), .Q(n191) );
  OAI212 U219 ( .A(n197), .B(n742), .C(n198), .Q(n196) );
  OAI212 U233 ( .A(n208), .B(n742), .C(n209), .Q(n207) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n742), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n791), .B(n742), .C(n789), .Q(n232) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U392 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U350 ( .A(n40), .B(n737), .C(n41), .Q(n39) );
  OAI212 U351 ( .A(n51), .B(n737), .C(n52), .Q(n50) );
  OAI212 U352 ( .A(n62), .B(n737), .C(n63), .Q(n61) );
  OAI212 U353 ( .A(n71), .B(n737), .C(n72), .Q(n70) );
  OAI212 U354 ( .A(n82), .B(n737), .C(n83), .Q(n81) );
  OAI212 U355 ( .A(n91), .B(n737), .C(n92), .Q(n90) );
  OAI212 U356 ( .A(n102), .B(n737), .C(n103), .Q(n101) );
  OAI212 U357 ( .A(n760), .B(n737), .C(n761), .Q(n108) );
  OAI212 U372 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U375 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NOR20 U349 ( .A(n205), .B(n212), .Q(n199) );
  BUF6 U358 ( .A(n2), .Q(n737) );
  OAI211 U359 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U360 ( .A(n245), .B(n241), .C(n242), .Q(n236) );
  AOI211 U361 ( .A(n200), .B(n183), .C(n184), .Q(n182) );
  NAND21 U362 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NOR21 U363 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND20 U364 ( .A(n780), .B(n206), .Q(n23) );
  NAND20 U365 ( .A(n778), .B(n195), .Q(n22) );
  NAND21 U366 ( .A(n790), .B(n242), .Q(n27) );
  NAND20 U367 ( .A(n782), .B(n213), .Q(n24) );
  INV0 U368 ( .A(n215), .Q(n786) );
  INV1 U369 ( .A(n247), .Q(n742) );
  INV0 U370 ( .A(n235), .Q(n791) );
  OAI210 U371 ( .A(n215), .B(n742), .C(n216), .Q(n214) );
  AOI210 U373 ( .A(n784), .B(n199), .C(n200), .Q(n198) );
  NAND20 U374 ( .A(n786), .B(n199), .Q(n197) );
  INV0 U376 ( .A(n216), .Q(n784) );
  INV0 U377 ( .A(n268), .Q(n741) );
  INV0 U378 ( .A(n199), .Q(n781) );
  OAI210 U379 ( .A(n176), .B(n737), .C(n177), .Q(n175) );
  OAI210 U380 ( .A(n213), .B(n205), .C(n206), .Q(n200) );
  OAI211 U381 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  OAI210 U382 ( .A(n244), .B(n742), .C(n245), .Q(n243) );
  NAND20 U383 ( .A(n235), .B(n787), .Q(n226) );
  AOI210 U384 ( .A(n236), .B(n787), .C(n788), .Q(n227) );
  NOR20 U385 ( .A(n192), .B(n781), .Q(n190) );
  OAI210 U386 ( .A(n274), .B(n740), .C(n275), .Q(n273) );
  INV0 U387 ( .A(n192), .Q(n778) );
  INV0 U388 ( .A(n271), .Q(n798) );
  INV1 U389 ( .A(n274), .Q(n799) );
  INV1 U390 ( .A(n252), .Q(n793) );
  INV0 U391 ( .A(n244), .Q(n792) );
  INV0 U393 ( .A(n241), .Q(n790) );
  INV0 U394 ( .A(n223), .Q(n785) );
  INV0 U395 ( .A(n205), .Q(n780) );
  INV0 U396 ( .A(n185), .Q(n777) );
  NOR20 U397 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NOR20 U398 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR20 U399 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NAND21 U400 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND21 U401 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NAND21 U402 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND21 U403 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND21 U404 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NAND20 U405 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NAND20 U406 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NAND20 U407 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND20 U408 ( .A(A[9]), .B(B[9]), .Q(n242) );
  NAND20 U409 ( .A(A[11]), .B(B[11]), .Q(n224) );
  NAND20 U410 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NAND20 U411 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NAND21 U412 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND20 U413 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NOR20 U414 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NOR21 U415 ( .A(n113), .B(n147), .Q(n4) );
  INV3 U416 ( .A(n147), .Q(n769) );
  NAND22 U417 ( .A(n4), .B(n42), .Q(n40) );
  AOI211 U418 ( .A(n3), .B(n42), .C(n43), .Q(n41) );
  NOR21 U419 ( .A(n44), .B(n75), .Q(n42) );
  NAND22 U420 ( .A(n4), .B(n53), .Q(n51) );
  AOI211 U421 ( .A(n3), .B(n53), .C(n54), .Q(n52) );
  NOR21 U422 ( .A(n747), .B(n75), .Q(n53) );
  NAND22 U423 ( .A(n4), .B(n93), .Q(n91) );
  AOI211 U424 ( .A(n3), .B(n93), .C(n94), .Q(n92) );
  NAND22 U425 ( .A(n4), .B(n751), .Q(n71) );
  AOI211 U426 ( .A(n3), .B(n751), .C(n752), .Q(n72) );
  INV3 U427 ( .A(n75), .Q(n751) );
  INV3 U428 ( .A(n167), .Q(n774) );
  INV3 U429 ( .A(n168), .Q(n775) );
  NAND22 U430 ( .A(n769), .B(n131), .Q(n129) );
  AOI211 U431 ( .A(n770), .B(n131), .C(n132), .Q(n130) );
  INV3 U432 ( .A(n4), .Q(n760) );
  INV3 U433 ( .A(n3), .Q(n761) );
  AOI211 U434 ( .A(n247), .B(n179), .C(n180), .Q(n2) );
  NOR21 U435 ( .A(n181), .B(n215), .Q(n179) );
  AOI211 U436 ( .A(n741), .B(n258), .C(n259), .Q(n257) );
  INV3 U437 ( .A(n236), .Q(n789) );
  NAND22 U438 ( .A(n93), .B(n77), .Q(n75) );
  INV3 U439 ( .A(n58), .Q(n748) );
  NAND22 U440 ( .A(n167), .B(n153), .Q(n147) );
  NAND22 U441 ( .A(n235), .B(n221), .Q(n215) );
  NAND22 U442 ( .A(n199), .B(n183), .Q(n181) );
  NAND22 U443 ( .A(n131), .B(n115), .Q(n113) );
  INV3 U444 ( .A(n148), .Q(n770) );
  INV3 U445 ( .A(n76), .Q(n752) );
  INV3 U446 ( .A(n131), .Q(n764) );
  INV3 U447 ( .A(n93), .Q(n755) );
  INV3 U448 ( .A(n57), .Q(n747) );
  INV3 U449 ( .A(n277), .Q(n740) );
  AOI211 U450 ( .A(n132), .B(n115), .C(n116), .Q(n114) );
  AOI211 U451 ( .A(n168), .B(n153), .C(n154), .Q(n148) );
  AOI211 U452 ( .A(n236), .B(n221), .C(n222), .Q(n216) );
  NAND22 U453 ( .A(n258), .B(n250), .Q(n248) );
  AOI211 U454 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR21 U455 ( .A(n252), .B(n255), .Q(n250) );
  NAND22 U456 ( .A(n4), .B(n757), .Q(n102) );
  AOI211 U457 ( .A(n3), .B(n757), .C(n758), .Q(n103) );
  INV3 U458 ( .A(n107), .Q(n758) );
  NAND22 U459 ( .A(n4), .B(n84), .Q(n82) );
  AOI211 U460 ( .A(n3), .B(n84), .C(n85), .Q(n83) );
  NOR21 U461 ( .A(n86), .B(n755), .Q(n84) );
  NAND22 U462 ( .A(n4), .B(n64), .Q(n62) );
  AOI211 U463 ( .A(n3), .B(n64), .C(n65), .Q(n63) );
  NOR21 U464 ( .A(n66), .B(n75), .Q(n64) );
  NAND22 U465 ( .A(n167), .B(n771), .Q(n158) );
  AOI211 U466 ( .A(n168), .B(n771), .C(n772), .Q(n159) );
  INV3 U467 ( .A(n163), .Q(n772) );
  NAND22 U468 ( .A(n769), .B(n766), .Q(n140) );
  AOI211 U469 ( .A(n770), .B(n766), .C(n767), .Q(n141) );
  INV3 U470 ( .A(n145), .Q(n767) );
  NAND22 U471 ( .A(n769), .B(n122), .Q(n120) );
  AOI211 U472 ( .A(n770), .B(n122), .C(n123), .Q(n121) );
  NOR21 U473 ( .A(n124), .B(n764), .Q(n122) );
  NOR21 U474 ( .A(n155), .B(n162), .Q(n153) );
  AOI211 U475 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U476 ( .A(n271), .B(n274), .Q(n269) );
  AOI211 U477 ( .A(n94), .B(n77), .C(n78), .Q(n76) );
  NOR21 U478 ( .A(n137), .B(n144), .Q(n131) );
  NOR21 U479 ( .A(n99), .B(n106), .Q(n93) );
  NOR21 U480 ( .A(n173), .B(n176), .Q(n167) );
  NOR21 U481 ( .A(n241), .B(n244), .Q(n235) );
  NOR21 U482 ( .A(n59), .B(n66), .Q(n57) );
  INV3 U483 ( .A(n231), .Q(n788) );
  NAND22 U484 ( .A(n786), .B(n782), .Q(n208) );
  AOI211 U485 ( .A(n784), .B(n782), .C(n783), .Q(n209) );
  INV3 U486 ( .A(n213), .Q(n783) );
  NAND22 U487 ( .A(n786), .B(n190), .Q(n188) );
  AOI211 U488 ( .A(n784), .B(n190), .C(n191), .Q(n189) );
  AOI211 U489 ( .A(n58), .B(n745), .C(n744), .Q(n45) );
  INV3 U490 ( .A(n49), .Q(n744) );
  NOR21 U491 ( .A(n185), .B(n192), .Q(n183) );
  NOR21 U492 ( .A(n79), .B(n86), .Q(n77) );
  NOR21 U493 ( .A(n117), .B(n124), .Q(n115) );
  AOI211 U494 ( .A(n741), .B(n796), .C(n797), .Q(n262) );
  INV3 U495 ( .A(n266), .Q(n797) );
  NOR21 U496 ( .A(n223), .B(n230), .Q(n221) );
  INV3 U497 ( .A(n132), .Q(n765) );
  NOR21 U498 ( .A(n260), .B(n265), .Q(n258) );
  NAND22 U499 ( .A(n57), .B(n745), .Q(n44) );
  INV3 U500 ( .A(n94), .Q(n756) );
  INV3 U501 ( .A(n200), .Q(n779) );
  INV3 U502 ( .A(n144), .Q(n766) );
  INV3 U503 ( .A(n106), .Q(n757) );
  INV3 U504 ( .A(n230), .Q(n787) );
  INV3 U505 ( .A(n212), .Q(n782) );
  INV3 U506 ( .A(n162), .Q(n771) );
  INV3 U507 ( .A(n265), .Q(n796) );
  INV3 U508 ( .A(n86), .Q(n753) );
  INV3 U509 ( .A(n66), .Q(n749) );
  INV3 U510 ( .A(n124), .Q(n762) );
  INV3 U511 ( .A(n155), .Q(n768) );
  INV3 U512 ( .A(n137), .Q(n763) );
  INV3 U513 ( .A(n117), .Q(n759) );
  INV3 U514 ( .A(n99), .Q(n754) );
  INV3 U515 ( .A(n79), .Q(n750) );
  INV3 U516 ( .A(n59), .Q(n746) );
  INV3 U517 ( .A(n176), .Q(n776) );
  INV3 U518 ( .A(n260), .Q(n795) );
  INV3 U519 ( .A(n173), .Q(n773) );
  INV3 U520 ( .A(n255), .Q(n794) );
  INV3 U521 ( .A(n278), .Q(n800) );
  NOR21 U522 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR21 U523 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NOR21 U524 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U525 ( .A(B[9]), .B(A[9]), .Q(n241) );
  NOR21 U526 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND22 U527 ( .A(A[17]), .B(B[17]), .Q(n174) );
  XNR21 U528 ( .A(n19), .B(n175), .Q(SUM[17]) );
  NAND22 U529 ( .A(n773), .B(n174), .Q(n19) );
  XNR21 U530 ( .A(n5), .B(n39), .Q(SUM[31]) );
  NAND22 U531 ( .A(n743), .B(n38), .Q(n5) );
  XNR21 U532 ( .A(n6), .B(n50), .Q(SUM[30]) );
  NAND22 U533 ( .A(n745), .B(n49), .Q(n6) );
  XNR21 U534 ( .A(n18), .B(n164), .Q(SUM[18]) );
  NAND22 U535 ( .A(n771), .B(n163), .Q(n18) );
  XNR21 U536 ( .A(n17), .B(n157), .Q(SUM[19]) );
  NAND22 U537 ( .A(n768), .B(n156), .Q(n17) );
  XNR21 U538 ( .A(n16), .B(n146), .Q(SUM[20]) );
  NAND22 U539 ( .A(n766), .B(n145), .Q(n16) );
  XNR21 U540 ( .A(n15), .B(n139), .Q(SUM[21]) );
  NAND22 U541 ( .A(n763), .B(n138), .Q(n15) );
  XNR21 U542 ( .A(n14), .B(n128), .Q(SUM[22]) );
  NAND22 U543 ( .A(n762), .B(n127), .Q(n14) );
  XNR21 U544 ( .A(n13), .B(n119), .Q(SUM[23]) );
  NAND22 U545 ( .A(n759), .B(n118), .Q(n13) );
  XNR21 U546 ( .A(n12), .B(n108), .Q(SUM[24]) );
  NAND22 U547 ( .A(n757), .B(n107), .Q(n12) );
  XNR21 U548 ( .A(n11), .B(n101), .Q(SUM[25]) );
  NAND22 U549 ( .A(n754), .B(n100), .Q(n11) );
  XNR21 U550 ( .A(n10), .B(n90), .Q(SUM[26]) );
  NAND22 U551 ( .A(n753), .B(n89), .Q(n10) );
  XNR21 U552 ( .A(n9), .B(n81), .Q(SUM[27]) );
  NAND22 U553 ( .A(n750), .B(n80), .Q(n9) );
  XNR21 U554 ( .A(n8), .B(n70), .Q(SUM[28]) );
  NAND22 U555 ( .A(n749), .B(n69), .Q(n8) );
  XNR21 U556 ( .A(n7), .B(n61), .Q(SUM[29]) );
  NAND22 U557 ( .A(n746), .B(n60), .Q(n7) );
  NOR21 U558 ( .A(B[22]), .B(A[22]), .Q(n124) );
  NOR21 U559 ( .A(B[26]), .B(A[26]), .Q(n86) );
  NOR21 U560 ( .A(B[28]), .B(A[28]), .Q(n66) );
  NOR21 U561 ( .A(B[14]), .B(A[14]), .Q(n192) );
  NOR21 U562 ( .A(B[29]), .B(A[29]), .Q(n59) );
  NOR21 U563 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR21 U564 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR21 U565 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR21 U566 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR21 U567 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR21 U568 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NOR21 U569 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR21 U570 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NOR21 U571 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U572 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NOR21 U573 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR21 U574 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR21 U575 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NOR21 U576 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND22 U577 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND22 U578 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NAND22 U579 ( .A(A[18]), .B(B[18]), .Q(n163) );
  XOR21 U580 ( .A(n28), .B(n742), .Q(SUM[8]) );
  NAND22 U581 ( .A(n792), .B(n245), .Q(n28) );
  XOR21 U582 ( .A(n20), .B(n737), .Q(SUM[16]) );
  NAND22 U583 ( .A(n776), .B(n177), .Q(n20) );
  XOR21 U584 ( .A(n30), .B(n257), .Q(SUM[6]) );
  NAND22 U585 ( .A(n794), .B(n256), .Q(n30) );
  NAND22 U586 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NAND22 U587 ( .A(A[28]), .B(B[28]), .Q(n69) );
  NAND22 U588 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NAND22 U589 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND22 U590 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NAND22 U591 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND22 U592 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND22 U593 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND22 U594 ( .A(A[29]), .B(B[29]), .Q(n60) );
  NAND22 U595 ( .A(A[5]), .B(B[5]), .Q(n261) );
  INV3 U596 ( .A(n48), .Q(n745) );
  NOR21 U597 ( .A(B[30]), .B(A[30]), .Q(n48) );
  XOR21 U598 ( .A(n31), .B(n262), .Q(SUM[5]) );
  NAND22 U599 ( .A(n795), .B(n261), .Q(n31) );
  XNR21 U600 ( .A(n29), .B(n254), .Q(SUM[7]) );
  NAND22 U601 ( .A(n793), .B(n253), .Q(n29) );
  XNR21 U602 ( .A(n27), .B(n243), .Q(SUM[9]) );
  XNR21 U603 ( .A(n26), .B(n232), .Q(SUM[10]) );
  NAND22 U604 ( .A(n787), .B(n231), .Q(n26) );
  XNR21 U605 ( .A(n25), .B(n225), .Q(SUM[11]) );
  NAND22 U606 ( .A(n785), .B(n224), .Q(n25) );
  XNR21 U607 ( .A(n24), .B(n214), .Q(SUM[12]) );
  XNR21 U608 ( .A(n23), .B(n207), .Q(SUM[13]) );
  XNR21 U609 ( .A(n22), .B(n196), .Q(SUM[14]) );
  XNR21 U610 ( .A(n21), .B(n187), .Q(SUM[15]) );
  NAND22 U611 ( .A(n777), .B(n186), .Q(n21) );
  XNR21 U612 ( .A(n32), .B(n741), .Q(SUM[4]) );
  NAND22 U613 ( .A(n796), .B(n266), .Q(n32) );
  NAND22 U614 ( .A(A[30]), .B(B[30]), .Q(n49) );
  INV3 U615 ( .A(n37), .Q(n743) );
  NOR21 U616 ( .A(A[31]), .B(B[31]), .Q(n37) );
  NAND22 U617 ( .A(B[31]), .B(A[31]), .Q(n38) );
  XOR21 U618 ( .A(n34), .B(n740), .Q(SUM[2]) );
  NAND22 U619 ( .A(n799), .B(n275), .Q(n34) );
  INV3 U620 ( .A(n280), .Q(n739) );
  NOR20 U621 ( .A(B[0]), .B(A[0]), .Q(n280) );
  INV3 U622 ( .A(n36), .Q(SUM[0]) );
  NAND22 U623 ( .A(n739), .B(n281), .Q(n36) );
  XNR21 U624 ( .A(n33), .B(n273), .Q(SUM[3]) );
  NAND22 U625 ( .A(n798), .B(n272), .Q(n33) );
  XOR21 U626 ( .A(n281), .B(n35), .Q(SUM[1]) );
  NAND22 U627 ( .A(n800), .B(n279), .Q(n35) );
  NAND20 U628 ( .A(A[0]), .B(B[0]), .Q(n281) );
endmodule


module adder_6 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_6_DW01_add_0 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n83, n84,
         n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n126, n127, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n141, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n422, n428, n434,
         n438, n440, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U91 ( .A(n521), .B(n102), .C(n103), .Q(n101) );
  OAI212 U105 ( .A(n152), .B(n113), .C(n114), .Q(n112) );
  OAI212 U165 ( .A(n158), .B(n521), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n580), .B(n521), .C(n578), .Q(n164) );
  AOI212 U195 ( .A(n179), .B(n247), .C(n180), .Q(n178) );
  OAI212 U197 ( .A(n181), .B(n220), .C(n182), .Q(n180) );
  OAI212 U207 ( .A(n188), .B(n526), .C(n189), .Q(n187) );
  OAI212 U219 ( .A(n197), .B(n526), .C(n198), .Q(n196) );
  OAI212 U233 ( .A(n208), .B(n526), .C(n209), .Q(n207) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n526), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n547), .B(n526), .C(n545), .Q(n232) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  OAI212 U306 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  OAI212 U323 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U329 ( .A(n274), .B(n524), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U492 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  OAI212 U499 ( .A(n173), .B(n177), .C(n174), .Q(n172) );
  OAI212 U512 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  AOI212 U381 ( .A(n153), .B(n172), .C(n154), .Q(n152) );
  OAI212 U427 ( .A(n252), .B(n256), .C(n253), .Q(n251) );
  OAI212 U459 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  OAI212 U464 ( .A(n120), .B(n521), .C(n121), .Q(n119) );
  OAI212 U495 ( .A(n573), .B(n521), .C(n570), .Q(n108) );
  OAI212 U514 ( .A(n42), .B(n521), .C(n43), .Q(n41) );
  OAI212 U533 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  OAI212 U540 ( .A(n155), .B(n163), .C(n156), .Q(n154) );
  OAI212 U511 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  NOR24 U349 ( .A(n223), .B(n230), .Q(n221) );
  OAI212 U350 ( .A(n88), .B(n564), .C(n89), .Q(n85) );
  NOR24 U351 ( .A(A[9]), .B(B[9]), .Q(n241) );
  INV10 U352 ( .A(n521), .Q(n527) );
  NOR22 U353 ( .A(A[5]), .B(B[5]), .Q(n260) );
  INV1 U354 ( .A(n244), .Q(n548) );
  NAND28 U355 ( .A(n550), .B(n537), .Q(n434) );
  NOR24 U356 ( .A(A[11]), .B(B[11]), .Q(n223) );
  NAND26 U357 ( .A(n171), .B(n153), .Q(n151) );
  AOI211 U358 ( .A(n520), .B(n97), .C(n98), .Q(n92) );
  OAI211 U359 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  AOI212 U360 ( .A(n520), .B(n66), .C(n67), .Q(n65) );
  NOR22 U361 ( .A(n70), .B(n6), .Q(n66) );
  NAND24 U362 ( .A(n65), .B(n438), .Q(n63) );
  CLKIN1 U363 ( .A(n536), .Q(n507) );
  NAND23 U364 ( .A(n557), .B(n527), .Q(n438) );
  NAND22 U365 ( .A(n111), .B(n97), .Q(n91) );
  NAND28 U366 ( .A(n97), .B(n77), .Q(n6) );
  NOR23 U367 ( .A(n99), .B(n106), .Q(n97) );
  NOR23 U368 ( .A(n117), .B(n126), .Q(n115) );
  NAND26 U369 ( .A(n434), .B(n206), .Q(n204) );
  NOR23 U370 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR22 U371 ( .A(B[8]), .B(A[8]), .Q(n244) );
  NOR23 U372 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NOR22 U373 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND22 U374 ( .A(A[29]), .B(B[29]), .Q(n62) );
  NAND22 U375 ( .A(B[8]), .B(A[8]), .Q(n245) );
  NAND22 U376 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U377 ( .A(A[10]), .B(B[10]), .Q(n231) );
  XNR21 U378 ( .A(n18), .B(n146), .Q(SUM[20]) );
  INV2 U379 ( .A(n97), .Q(n566) );
  INV2 U380 ( .A(n219), .Q(n541) );
  NOR23 U382 ( .A(n181), .B(n219), .Q(n179) );
  OAI211 U383 ( .A(n129), .B(n521), .C(n130), .Q(n128) );
  NOR21 U384 ( .A(n126), .B(n577), .Q(n122) );
  INV3 U385 ( .A(n542), .Q(n504) );
  NOR23 U386 ( .A(n162), .B(n155), .Q(n153) );
  NAND24 U387 ( .A(n518), .B(n111), .Q(n428) );
  BUF2 U388 ( .A(n137), .Q(n505) );
  AOI212 U389 ( .A(n60), .B(n560), .C(n559), .Q(n47) );
  NAND26 U390 ( .A(n203), .B(n183), .Q(n181) );
  NAND21 U391 ( .A(B[23]), .B(A[23]), .Q(n118) );
  NOR23 U392 ( .A(A[27]), .B(B[27]), .Q(n79) );
  NOR23 U393 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NAND22 U394 ( .A(B[24]), .B(A[24]), .Q(n107) );
  CLKIN3 U395 ( .A(n144), .Q(n584) );
  NAND20 U396 ( .A(n584), .B(n145), .Q(n18) );
  INV0 U397 ( .A(n145), .Q(n585) );
  CLKIN0 U398 ( .A(n163), .Q(n568) );
  INV1 U399 ( .A(n60), .Q(n552) );
  NOR23 U400 ( .A(n61), .B(n70), .Q(n59) );
  NAND23 U401 ( .A(n440), .B(n54), .Q(n52) );
  INV1 U402 ( .A(n162), .Q(n571) );
  INV0 U403 ( .A(n505), .Q(n576) );
  CLKIN1 U404 ( .A(n575), .Q(n508) );
  NAND21 U405 ( .A(n560), .B(n51), .Q(n8) );
  NAND22 U406 ( .A(B[19]), .B(A[19]), .Q(n156) );
  NAND21 U407 ( .A(n582), .B(n107), .Q(n14) );
  INV1 U408 ( .A(n107), .Q(n581) );
  NAND22 U409 ( .A(n111), .B(n66), .Q(n64) );
  NAND26 U410 ( .A(n135), .B(n115), .Q(n113) );
  INV2 U411 ( .A(n135), .Q(n577) );
  NOR24 U412 ( .A(n137), .B(n144), .Q(n135) );
  NAND21 U413 ( .A(n111), .B(n582), .Q(n102) );
  NAND21 U414 ( .A(n111), .B(n563), .Q(n73) );
  NAND22 U415 ( .A(n111), .B(n55), .Q(n53) );
  NAND22 U416 ( .A(B[25]), .B(A[25]), .Q(n100) );
  AOI211 U417 ( .A(n520), .B(n44), .C(n45), .Q(n43) );
  OAI212 U418 ( .A(n5), .B(n46), .C(n47), .Q(n45) );
  NAND23 U419 ( .A(B[14]), .B(A[14]), .Q(n195) );
  NAND22 U420 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NOR24 U421 ( .A(B[15]), .B(A[15]), .Q(n511) );
  AOI211 U422 ( .A(n569), .B(n135), .C(n508), .Q(n130) );
  INV1 U423 ( .A(n569), .Q(n513) );
  NAND22 U424 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NAND21 U425 ( .A(n565), .B(n100), .Q(n13) );
  CLKIN3 U426 ( .A(n247), .Q(n526) );
  BUF2 U428 ( .A(n194), .Q(n506) );
  NAND20 U429 ( .A(n239), .B(n543), .Q(n226) );
  INV1 U430 ( .A(n204), .Q(n536) );
  NAND24 U431 ( .A(A[12]), .B(B[12]), .Q(n213) );
  INV2 U432 ( .A(n136), .Q(n575) );
  BUF2 U433 ( .A(n259), .Q(n509) );
  INV3 U434 ( .A(n6), .Q(n563) );
  INV1 U435 ( .A(n126), .Q(n587) );
  NOR24 U436 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NAND22 U437 ( .A(n92), .B(n422), .Q(n90) );
  INV0 U438 ( .A(n550), .Q(n510) );
  NOR23 U439 ( .A(n205), .B(n212), .Q(n203) );
  NAND23 U440 ( .A(B[16]), .B(A[16]), .Q(n177) );
  OAI211 U441 ( .A(n140), .B(n521), .C(n141), .Q(n139) );
  AOI211 U442 ( .A(n569), .B(n584), .C(n585), .Q(n141) );
  CLKIN3 U443 ( .A(n61), .Q(n553) );
  NAND22 U444 ( .A(A[21]), .B(B[21]), .Q(n138) );
  INV4 U445 ( .A(n517), .Q(n518) );
  INV0 U446 ( .A(n79), .Q(n583) );
  NAND22 U447 ( .A(A[13]), .B(B[13]), .Q(n206) );
  INV6 U448 ( .A(n213), .Q(n550) );
  NAND21 U449 ( .A(n258), .B(n250), .Q(n248) );
  XNR22 U450 ( .A(n15), .B(n119), .Q(SUM[23]) );
  XNR22 U451 ( .A(n52), .B(n8), .Q(SUM[30]) );
  NAND21 U452 ( .A(A[27]), .B(B[27]), .Q(n80) );
  INV2 U453 ( .A(n98), .Q(n564) );
  AOI210 U454 ( .A(n569), .B(n122), .C(n123), .Q(n121) );
  NAND24 U455 ( .A(n428), .B(n83), .Q(n81) );
  CLKIN15 U456 ( .A(n519), .Q(n520) );
  NAND22 U457 ( .A(A[28]), .B(B[28]), .Q(n71) );
  INV0 U458 ( .A(n155), .Q(n574) );
  BUF15 U460 ( .A(n178), .Q(n521) );
  INV0 U461 ( .A(n99), .Q(n565) );
  NOR24 U462 ( .A(B[25]), .B(A[25]), .Q(n99) );
  XNR22 U463 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI211 U465 ( .A(n151), .B(n521), .C(n513), .Q(n146) );
  INV6 U466 ( .A(n112), .Q(n519) );
  XNR22 U467 ( .A(n9), .B(n63), .Q(SUM[29]) );
  NOR23 U468 ( .A(n46), .B(n6), .Q(n44) );
  NAND24 U469 ( .A(n59), .B(n560), .Q(n46) );
  NOR23 U470 ( .A(n555), .B(n6), .Q(n55) );
  CLKIN6 U471 ( .A(n59), .Q(n555) );
  OAI211 U472 ( .A(n176), .B(n521), .C(n177), .Q(n175) );
  NOR24 U473 ( .A(n79), .B(n88), .Q(n77) );
  XNR22 U474 ( .A(n13), .B(n101), .Q(SUM[25]) );
  INV0 U475 ( .A(n176), .Q(n586) );
  OAI211 U476 ( .A(n126), .B(n575), .C(n127), .Q(n123) );
  OAI210 U477 ( .A(n177), .B(n173), .C(n174), .Q(n516) );
  NOR22 U478 ( .A(n173), .B(n176), .Q(n171) );
  NOR23 U479 ( .A(A[18]), .B(B[18]), .Q(n162) );
  INV0 U480 ( .A(n173), .Q(n579) );
  XNR22 U481 ( .A(n7), .B(n41), .Q(SUM[31]) );
  INV2 U482 ( .A(n223), .Q(n540) );
  BUF2 U483 ( .A(n511), .Q(n512) );
  INV0 U484 ( .A(n512), .Q(n539) );
  AOI212 U485 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  AOI212 U486 ( .A(n520), .B(n55), .C(n56), .Q(n54) );
  INV2 U487 ( .A(n152), .Q(n569) );
  BUF2 U488 ( .A(n194), .Q(n514) );
  NAND21 U489 ( .A(n171), .B(n571), .Q(n158) );
  INV1 U490 ( .A(n171), .Q(n580) );
  INV2 U491 ( .A(n111), .Q(n573) );
  NAND22 U493 ( .A(A[26]), .B(B[26]), .Q(n89) );
  INV0 U494 ( .A(n514), .Q(n549) );
  NAND22 U496 ( .A(B[9]), .B(A[9]), .Q(n242) );
  NOR24 U497 ( .A(B[21]), .B(A[21]), .Q(n137) );
  INV0 U498 ( .A(n241), .Q(n546) );
  NAND21 U500 ( .A(n572), .B(n584), .Q(n140) );
  INV2 U501 ( .A(n151), .Q(n572) );
  NAND22 U502 ( .A(B[17]), .B(A[17]), .Q(n174) );
  NOR24 U503 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR20 U504 ( .A(n506), .B(n538), .Q(n190) );
  NOR24 U505 ( .A(A[19]), .B(B[19]), .Q(n155) );
  XNR22 U506 ( .A(n10), .B(n72), .Q(SUM[28]) );
  OAI212 U507 ( .A(n73), .B(n521), .C(n74), .Q(n72) );
  BUF2 U508 ( .A(n240), .Q(n515) );
  OAI210 U509 ( .A(n514), .B(n536), .C(n195), .Q(n191) );
  INV1 U510 ( .A(n220), .Q(n542) );
  INV0 U513 ( .A(n252), .Q(n532) );
  INV2 U515 ( .A(n5), .Q(n561) );
  OAI212 U516 ( .A(n5), .B(n555), .C(n552), .Q(n56) );
  INV6 U517 ( .A(n205), .Q(n537) );
  NOR24 U518 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NOR24 U519 ( .A(n241), .B(n244), .Q(n239) );
  NAND22 U520 ( .A(B[18]), .B(A[18]), .Q(n163) );
  OAI212 U521 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  NOR23 U522 ( .A(A[26]), .B(B[26]), .Q(n88) );
  NOR24 U523 ( .A(B[23]), .B(A[23]), .Q(n117) );
  INV3 U524 ( .A(n106), .Q(n582) );
  XNR22 U525 ( .A(n11), .B(n81), .Q(SUM[27]) );
  CLKIN2 U526 ( .A(n203), .Q(n538) );
  OAI212 U527 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  AOI212 U528 ( .A(n520), .B(n563), .C(n561), .Q(n74) );
  NOR24 U529 ( .A(A[17]), .B(B[17]), .Q(n173) );
  NAND21 U530 ( .A(n572), .B(n135), .Q(n129) );
  OAI211 U531 ( .A(n244), .B(n526), .C(n245), .Q(n243) );
  NOR24 U532 ( .A(A[14]), .B(B[14]), .Q(n194) );
  AOI212 U534 ( .A(n183), .B(n204), .C(n184), .Q(n182) );
  NAND21 U535 ( .A(B[11]), .B(A[11]), .Q(n224) );
  OAI212 U536 ( .A(n195), .B(n511), .C(n186), .Q(n184) );
  AOI211 U537 ( .A(n520), .B(n582), .C(n581), .Q(n103) );
  AOI211 U538 ( .A(n520), .B(n84), .C(n85), .Q(n83) );
  NOR24 U539 ( .A(n113), .B(n151), .Q(n111) );
  NAND21 U541 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND21 U542 ( .A(A[7]), .B(B[7]), .Q(n253) );
  AOI212 U543 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  NOR22 U544 ( .A(n252), .B(n255), .Q(n250) );
  NAND24 U545 ( .A(n221), .B(n239), .Q(n219) );
  OAI211 U546 ( .A(n219), .B(n526), .C(n504), .Q(n214) );
  NOR24 U547 ( .A(n185), .B(n194), .Q(n183) );
  NOR23 U548 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NOR24 U549 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND22 U550 ( .A(n549), .B(n195), .Q(n24) );
  NAND22 U551 ( .A(n84), .B(n527), .Q(n517) );
  NAND22 U552 ( .A(A[22]), .B(B[22]), .Q(n127) );
  CLKIN0 U553 ( .A(n515), .Q(n545) );
  CLKIN0 U554 ( .A(n516), .Q(n578) );
  NAND21 U555 ( .A(n572), .B(n122), .Q(n120) );
  NOR22 U556 ( .A(B[16]), .B(A[16]), .Q(n176) );
  INV0 U557 ( .A(n212), .Q(n551) );
  INV0 U558 ( .A(n266), .Q(n534) );
  NAND22 U559 ( .A(n527), .B(n567), .Q(n422) );
  AOI210 U560 ( .A(n542), .B(n203), .C(n507), .Q(n198) );
  NAND20 U561 ( .A(n541), .B(n203), .Q(n197) );
  CLKIN0 U562 ( .A(n239), .Q(n547) );
  AOI210 U563 ( .A(n525), .B(n258), .C(n509), .Q(n257) );
  INV0 U564 ( .A(n260), .Q(n533) );
  INV0 U565 ( .A(n230), .Q(n543) );
  NOR20 U566 ( .A(n260), .B(n265), .Q(n258) );
  NOR22 U567 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR22 U568 ( .A(B[6]), .B(A[6]), .Q(n255) );
  NAND21 U569 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND21 U570 ( .A(A[31]), .B(B[31]), .Q(n40) );
  INV2 U571 ( .A(n39), .Q(n558) );
  XOR21 U572 ( .A(n30), .B(n526), .Q(SUM[8]) );
  INV3 U573 ( .A(n53), .Q(n554) );
  INV3 U574 ( .A(n520), .Q(n570) );
  NAND20 U575 ( .A(n541), .B(n551), .Q(n208) );
  AOI210 U576 ( .A(n542), .B(n551), .C(n550), .Q(n209) );
  NAND22 U577 ( .A(n554), .B(n527), .Q(n440) );
  INV3 U578 ( .A(n91), .Q(n567) );
  INV3 U579 ( .A(n64), .Q(n557) );
  INV3 U580 ( .A(n268), .Q(n525) );
  NOR21 U581 ( .A(n88), .B(n566), .Q(n84) );
  INV3 U582 ( .A(n231), .Q(n544) );
  INV3 U583 ( .A(n51), .Q(n559) );
  NAND20 U584 ( .A(n541), .B(n190), .Q(n188) );
  AOI210 U585 ( .A(n542), .B(n190), .C(n191), .Q(n189) );
  NAND22 U586 ( .A(n533), .B(n261), .Q(n33) );
  INV3 U587 ( .A(n70), .Q(n556) );
  INV3 U588 ( .A(n255), .Q(n531) );
  NAND22 U589 ( .A(n529), .B(n272), .Q(n35) );
  INV3 U590 ( .A(n271), .Q(n529) );
  INV3 U591 ( .A(n278), .Q(n528) );
  INV3 U592 ( .A(n265), .Q(n535) );
  INV3 U593 ( .A(n274), .Q(n530) );
  AOI211 U594 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  NOR21 U595 ( .A(n271), .B(n274), .Q(n269) );
  INV3 U596 ( .A(n277), .Q(n524) );
  NOR21 U597 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR21 U598 ( .A(B[1]), .B(A[1]), .Q(n278) );
  INV3 U599 ( .A(n50), .Q(n560) );
  NOR21 U600 ( .A(B[30]), .B(A[30]), .Q(n50) );
  NOR21 U601 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NOR21 U602 ( .A(B[4]), .B(A[4]), .Q(n265) );
  NAND22 U603 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND22 U604 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND22 U605 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NOR21 U606 ( .A(B[31]), .B(A[31]), .Q(n39) );
  INV3 U607 ( .A(n280), .Q(n523) );
  NOR21 U608 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND22 U609 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U610 ( .A(n553), .B(n62), .Q(n9) );
  NAND22 U611 ( .A(n558), .B(n40), .Q(n7) );
  NAND20 U612 ( .A(n562), .B(n89), .Q(n12) );
  XNR21 U613 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND20 U614 ( .A(n587), .B(n127), .Q(n16) );
  NAND20 U615 ( .A(n556), .B(n71), .Q(n10) );
  XOR20 U616 ( .A(n22), .B(n521), .Q(SUM[16]) );
  NAND20 U617 ( .A(n586), .B(n177), .Q(n22) );
  XNR21 U618 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND20 U619 ( .A(n537), .B(n206), .Q(n25) );
  XNR21 U620 ( .A(n23), .B(n187), .Q(SUM[15]) );
  NAND20 U621 ( .A(n186), .B(n539), .Q(n23) );
  XNR21 U622 ( .A(n29), .B(n243), .Q(SUM[9]) );
  NAND20 U623 ( .A(n546), .B(n242), .Q(n29) );
  XNR21 U624 ( .A(n26), .B(n214), .Q(SUM[12]) );
  NAND20 U625 ( .A(n551), .B(n510), .Q(n26) );
  XNR21 U626 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NAND20 U627 ( .A(n543), .B(n231), .Q(n28) );
  XNR21 U628 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND20 U629 ( .A(n583), .B(n80), .Q(n11) );
  XNR21 U630 ( .A(n24), .B(n196), .Q(SUM[14]) );
  XNR21 U631 ( .A(n27), .B(n225), .Q(SUM[11]) );
  NAND20 U632 ( .A(n540), .B(n224), .Q(n27) );
  NAND20 U633 ( .A(n548), .B(n245), .Q(n30) );
  XOR21 U634 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI211 U635 ( .A(n525), .B(n535), .C(n534), .Q(n262) );
  XOR21 U636 ( .A(n32), .B(n257), .Q(SUM[6]) );
  NAND20 U637 ( .A(n531), .B(n256), .Q(n32) );
  XNR21 U638 ( .A(n31), .B(n254), .Q(SUM[7]) );
  NAND20 U639 ( .A(n532), .B(n253), .Q(n31) );
  XNR21 U640 ( .A(n21), .B(n175), .Q(SUM[17]) );
  NAND20 U641 ( .A(n174), .B(n579), .Q(n21) );
  XNR21 U642 ( .A(n19), .B(n157), .Q(SUM[19]) );
  NAND20 U643 ( .A(n574), .B(n156), .Q(n19) );
  XNR21 U644 ( .A(n17), .B(n139), .Q(SUM[21]) );
  NAND20 U645 ( .A(n576), .B(n138), .Q(n17) );
  NAND20 U646 ( .A(n588), .B(n118), .Q(n15) );
  XNR21 U647 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR21 U648 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NAND20 U649 ( .A(n163), .B(n571), .Q(n20) );
  XOR21 U650 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U651 ( .A(n528), .B(n279), .Q(n37) );
  XNR21 U652 ( .A(n34), .B(n525), .Q(SUM[4]) );
  NAND20 U653 ( .A(n535), .B(n266), .Q(n34) );
  XOR21 U654 ( .A(n36), .B(n524), .Q(SUM[2]) );
  NAND22 U655 ( .A(n530), .B(n275), .Q(n36) );
  INV3 U656 ( .A(n38), .Q(SUM[0]) );
  NAND22 U657 ( .A(n523), .B(n281), .Q(n38) );
  NAND22 U658 ( .A(n111), .B(n44), .Q(n42) );
  CLKIN0 U659 ( .A(n88), .Q(n562) );
  NAND22 U660 ( .A(A[20]), .B(B[20]), .Q(n145) );
  INV2 U661 ( .A(n117), .Q(n588) );
  AOI210 U662 ( .A(n515), .B(n543), .C(n544), .Q(n227) );
  AOI210 U663 ( .A(n516), .B(n571), .C(n568), .Q(n159) );
endmodule


module adder_5 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_5_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n62, n67,
         n68, n69, n70, n71, n74, n75, n76, n81, n82, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n95, n96, n97, n98, n99, n100, n105, n106, n107,
         n108, n109, n112, n113, n114, n115, n116, n121, n122, n123, n124,
         n125, n126, n127, n130, n131, n132, n135, n136, n141, n142, n143,
         n144, n145, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n163, n164, n165, n166, n167, n168,
         n173, n174, n175, n176, n177, n180, n181, n182, n183, n184, n189,
         n190, n191, n192, n193, n194, n195, n198, n199, n200, n203, n204,
         n209, n210, n211, n212, n213, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n228, n229, n230, n231, n236, n237,
         n238, n241, n242, n244, n245, n246, n247, n248, n249, n250, n251,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n265, n266, n267, n268, n269, n405, n411, n419, n420, n556, n700,
         n703, n704, n707, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863;

  OAI212 U60 ( .A(n818), .B(n796), .C(n817), .Q(n76) );
  OAI212 U64 ( .A(n81), .B(n116), .C(n82), .Q(n2) );
  OAI212 U74 ( .A(n88), .B(n796), .C(n89), .Q(n87) );
  OAI212 U86 ( .A(n97), .B(n796), .C(n98), .Q(n96) );
  AOI212 U116 ( .A(n136), .B(n121), .C(n122), .Q(n116) );
  OAI212 U124 ( .A(n126), .B(n796), .C(n127), .Q(n125) );
  OAI212 U134 ( .A(n842), .B(n796), .C(n839), .Q(n132) );
  AOI212 U208 ( .A(n204), .B(n189), .C(n190), .Q(n184) );
  OAI212 U247 ( .A(n216), .B(n244), .C(n217), .Q(n215) );
  OAI212 U251 ( .A(n220), .B(n228), .C(n221), .Q(n219) );
  OAI212 U273 ( .A(n242), .B(n236), .C(n237), .Q(n231) );
  OAI212 U311 ( .A(n263), .B(n259), .C(n260), .Q(n258) );
  OAI212 U317 ( .A(n262), .B(n799), .C(n263), .Q(n261) );
  OAI212 U324 ( .A(n269), .B(n266), .C(n267), .Q(n265) );
  OAI212 U600 ( .A(n115), .B(n796), .C(n116), .Q(n114) );
  OAI212 U466 ( .A(n181), .B(n173), .C(n174), .Q(n168) );
  AOI212 U344 ( .A(n777), .B(n147), .C(n148), .Q(n1) );
  OAI212 U425 ( .A(n213), .B(n209), .C(n210), .Q(n204) );
  OAI212 U451 ( .A(n145), .B(n794), .C(n142), .Q(n136) );
  OAI212 U437 ( .A(n199), .B(n191), .C(n192), .Q(n190) );
  OAI212 U345 ( .A(n70), .B(n783), .C(n71), .Q(n69) );
  OAI212 U406 ( .A(n213), .B(n209), .C(n210), .Q(n405) );
  OAI212 U438 ( .A(n75), .B(n67), .C(n68), .Q(n62) );
  OAI212 U511 ( .A(n256), .B(n254), .C(n255), .Q(n253) );
  OAI212 U457 ( .A(n251), .B(n247), .C(n248), .Q(n246) );
  AOI212 U499 ( .A(n253), .B(n245), .C(n246), .Q(n244) );
  OAI212 U623 ( .A(n184), .B(n149), .C(n150), .Q(n148) );
  OAI212 U375 ( .A(n250), .B(n800), .C(n251), .Q(n249) );
  OAI212 U445 ( .A(n165), .B(n802), .C(n166), .Q(n164) );
  OAI212 U453 ( .A(n194), .B(n802), .C(n195), .Q(n193) );
  XNR22 U337 ( .A(n19), .B(n175), .Q(SUM[16]) );
  INV8 U338 ( .A(n777), .Q(n802) );
  NAND21 U339 ( .A(n825), .B(n158), .Q(n156) );
  NAND21 U340 ( .A(n824), .B(n777), .Q(n700) );
  NAND21 U341 ( .A(n849), .B(n248), .Q(n29) );
  AOI212 U342 ( .A(n2), .B(n52), .C(n53), .Q(n51) );
  NOR22 U343 ( .A(B[22]), .B(A[22]), .Q(n123) );
  NAND21 U346 ( .A(n203), .B(n777), .Q(n707) );
  INV12 U347 ( .A(n776), .Q(n777) );
  XOR22 U348 ( .A(n27), .B(n238), .Q(SUM[8]) );
  NAND24 U349 ( .A(n230), .B(n218), .Q(n216) );
  INV6 U350 ( .A(n802), .Q(n792) );
  NAND21 U351 ( .A(A[22]), .B(B[22]), .Q(n124) );
  NOR24 U352 ( .A(n220), .B(n225), .Q(n218) );
  NOR22 U353 ( .A(n794), .B(n144), .Q(n135) );
  NOR24 U354 ( .A(B[7]), .B(A[7]), .Q(n241) );
  NOR24 U355 ( .A(n241), .B(n236), .Q(n230) );
  NAND26 U356 ( .A(n836), .B(n803), .Q(n704) );
  BUF15 U357 ( .A(n1), .Q(n796) );
  NOR23 U358 ( .A(n209), .B(n212), .Q(n203) );
  NOR24 U359 ( .A(A[12]), .B(B[12]), .Q(n209) );
  NAND26 U360 ( .A(n703), .B(n704), .Q(SUM[13]) );
  NOR22 U361 ( .A(B[24]), .B(A[24]), .Q(n105) );
  XOR22 U362 ( .A(n26), .B(n229), .Q(SUM[9]) );
  INV6 U363 ( .A(n215), .Q(n776) );
  NOR22 U364 ( .A(B[13]), .B(A[13]), .Q(n198) );
  NAND23 U365 ( .A(n99), .B(n819), .Q(n81) );
  NOR21 U366 ( .A(B[25]), .B(A[25]), .Q(n92) );
  NAND24 U367 ( .A(n203), .B(n189), .Q(n183) );
  AOI211 U368 ( .A(n100), .B(n819), .C(n84), .Q(n82) );
  CLKIN3 U369 ( .A(n182), .Q(n789) );
  NOR22 U370 ( .A(n191), .B(n198), .Q(n189) );
  INV3 U371 ( .A(n92), .Q(n821) );
  NOR22 U372 ( .A(n795), .B(n130), .Q(n121) );
  NAND23 U373 ( .A(A[11]), .B(B[11]), .Q(n213) );
  INV3 U374 ( .A(n99), .Q(n852) );
  NOR21 U376 ( .A(B[20]), .B(A[20]), .Q(n141) );
  INV6 U377 ( .A(n782), .Q(n783) );
  INV3 U378 ( .A(n62), .Q(n814) );
  NAND23 U379 ( .A(n135), .B(n121), .Q(n115) );
  AOI211 U380 ( .A(n840), .B(n855), .C(n854), .Q(n109) );
  XOR21 U381 ( .A(n25), .B(n222), .Q(SUM[10]) );
  NAND23 U382 ( .A(n790), .B(n791), .Q(SUM[15]) );
  INV2 U383 ( .A(n231), .Q(n830) );
  NOR22 U384 ( .A(B[11]), .B(A[11]), .Q(n212) );
  NAND22 U385 ( .A(A[13]), .B(B[13]), .Q(n199) );
  INV3 U386 ( .A(n184), .Q(n822) );
  OAI211 U387 ( .A(n57), .B(n47), .C(n48), .Q(n46) );
  NOR21 U388 ( .A(n47), .B(n54), .Q(n45) );
  INV3 U389 ( .A(n822), .Q(n778) );
  INV3 U390 ( .A(n199), .Q(n838) );
  INV2 U391 ( .A(n830), .Q(n779) );
  INV3 U392 ( .A(n849), .Q(n780) );
  INV3 U393 ( .A(n116), .Q(n840) );
  AOI211 U394 ( .A(n2), .B(n815), .C(n62), .Q(n60) );
  AOI211 U395 ( .A(n2), .B(n816), .C(n813), .Q(n71) );
  NOR23 U396 ( .A(n173), .B(n180), .Q(n167) );
  CLKIN1 U397 ( .A(n230), .Q(n832) );
  BUF6 U398 ( .A(n228), .Q(n781) );
  CLKIN1 U399 ( .A(n247), .Q(n849) );
  NAND21 U400 ( .A(n96), .B(n10), .Q(n786) );
  CLKIN3 U401 ( .A(n96), .Q(n784) );
  CLKIN4 U402 ( .A(n796), .Q(n782) );
  NAND22 U403 ( .A(n784), .B(n785), .Q(n787) );
  NAND24 U404 ( .A(n786), .B(n787), .Q(SUM[25]) );
  INV2 U405 ( .A(n10), .Q(n785) );
  OAI210 U407 ( .A(n39), .B(n783), .C(n40), .Q(n38) );
  NAND21 U408 ( .A(n237), .B(n861), .Q(n27) );
  NAND24 U409 ( .A(A[7]), .B(B[7]), .Q(n242) );
  NAND23 U410 ( .A(B[8]), .B(A[8]), .Q(n237) );
  NAND22 U411 ( .A(A[9]), .B(B[9]), .Q(n228) );
  NAND22 U412 ( .A(n20), .B(n182), .Q(n790) );
  NAND22 U413 ( .A(n788), .B(n789), .Q(n791) );
  INV3 U414 ( .A(n20), .Q(n788) );
  NAND20 U415 ( .A(n857), .B(n181), .Q(n20) );
  INV1 U416 ( .A(n241), .Q(n831) );
  NOR20 U417 ( .A(n225), .B(n832), .Q(n223) );
  NOR24 U418 ( .A(B[9]), .B(A[9]), .Q(n225) );
  OAI212 U419 ( .A(n113), .B(n105), .C(n106), .Q(n100) );
  NAND21 U420 ( .A(A[23]), .B(B[23]), .Q(n113) );
  NAND24 U421 ( .A(n848), .B(n792), .Q(n793) );
  NAND28 U422 ( .A(n793), .B(n213), .Q(n211) );
  XNR22 U423 ( .A(n164), .B(n18), .Q(SUM[17]) );
  NOR21 U424 ( .A(B[26]), .B(A[26]), .Q(n85) );
  INV2 U426 ( .A(n115), .Q(n843) );
  NAND21 U427 ( .A(A[21]), .B(B[21]), .Q(n131) );
  NOR24 U428 ( .A(B[10]), .B(A[10]), .Q(n220) );
  NAND24 U429 ( .A(n167), .B(n151), .Q(n149) );
  NAND24 U430 ( .A(A[5]), .B(B[5]), .Q(n251) );
  OAI212 U431 ( .A(n163), .B(n153), .C(n154), .Q(n152) );
  NAND21 U432 ( .A(A[18]), .B(B[18]), .Q(n154) );
  NOR23 U433 ( .A(B[16]), .B(A[16]), .Q(n173) );
  NOR24 U434 ( .A(B[6]), .B(A[6]), .Q(n247) );
  NAND22 U435 ( .A(B[6]), .B(A[6]), .Q(n248) );
  CLKIN3 U436 ( .A(n160), .Q(n853) );
  OAI210 U439 ( .A(n160), .B(n835), .C(n163), .Q(n159) );
  NOR21 U440 ( .A(n160), .B(n834), .Q(n158) );
  NOR23 U441 ( .A(n153), .B(n160), .Q(n151) );
  NAND21 U442 ( .A(A[17]), .B(B[17]), .Q(n163) );
  NAND21 U443 ( .A(A[16]), .B(B[16]), .Q(n174) );
  NAND21 U444 ( .A(A[20]), .B(B[20]), .Q(n142) );
  NOR22 U446 ( .A(B[17]), .B(A[17]), .Q(n160) );
  NAND21 U447 ( .A(A[14]), .B(B[14]), .Q(n192) );
  OAI212 U448 ( .A(n131), .B(n795), .C(n124), .Q(n122) );
  INV2 U449 ( .A(n2), .Q(n817) );
  OAI212 U450 ( .A(n108), .B(n796), .C(n109), .Q(n107) );
  XNR22 U452 ( .A(n17), .B(n155), .Q(SUM[18]) );
  NAND22 U454 ( .A(n3), .B(n52), .Q(n50) );
  NOR21 U455 ( .A(n54), .B(n411), .Q(n52) );
  NOR24 U456 ( .A(B[8]), .B(A[8]), .Q(n236) );
  CLKIN6 U458 ( .A(n200), .Q(n803) );
  OAI212 U459 ( .A(n59), .B(n783), .C(n60), .Q(n58) );
  INV2 U460 ( .A(n225), .Q(n828) );
  OAI210 U461 ( .A(n225), .B(n830), .C(n781), .Q(n224) );
  XNR22 U462 ( .A(n6), .B(n58), .Q(SUM[29]) );
  NAND20 U463 ( .A(n816), .B(n75), .Q(n8) );
  NAND21 U464 ( .A(A[27]), .B(B[27]), .Q(n75) );
  NAND21 U465 ( .A(A[10]), .B(B[10]), .Q(n221) );
  INV0 U467 ( .A(n220), .Q(n827) );
  XNR21 U468 ( .A(n28), .B(n801), .Q(SUM[7]) );
  OAI211 U469 ( .A(n54), .B(n814), .C(n57), .Q(n53) );
  NOR21 U470 ( .A(B[29]), .B(A[29]), .Q(n54) );
  OAI211 U471 ( .A(n50), .B(n796), .C(n51), .Q(n49) );
  XOR22 U472 ( .A(n16), .B(n796), .Q(SUM[19]) );
  XNR22 U473 ( .A(n11), .B(n107), .Q(SUM[24]) );
  XNR22 U474 ( .A(n8), .B(n76), .Q(SUM[27]) );
  NOR22 U475 ( .A(B[15]), .B(A[15]), .Q(n180) );
  NAND22 U476 ( .A(A[15]), .B(B[15]), .Q(n181) );
  OAI212 U477 ( .A(n144), .B(n796), .C(n145), .Q(n143) );
  INV0 U478 ( .A(n236), .Q(n861) );
  INV2 U479 ( .A(n180), .Q(n857) );
  XNR22 U480 ( .A(n132), .B(n14), .Q(SUM[21]) );
  XNR22 U481 ( .A(n12), .B(n114), .Q(SUM[23]) );
  NAND20 U482 ( .A(n855), .B(n113), .Q(n12) );
  INV1 U483 ( .A(n113), .Q(n854) );
  XNR22 U484 ( .A(n23), .B(n211), .Q(SUM[12]) );
  XNR22 U485 ( .A(n13), .B(n125), .Q(SUM[22]) );
  OAI212 U486 ( .A(n183), .B(n802), .C(n778), .Q(n182) );
  XNR22 U487 ( .A(n15), .B(n143), .Q(SUM[20]) );
  NOR22 U488 ( .A(n105), .B(n112), .Q(n99) );
  NOR21 U489 ( .A(B[23]), .B(A[23]), .Q(n112) );
  AOI211 U490 ( .A(n840), .B(n99), .C(n100), .Q(n98) );
  NAND22 U491 ( .A(n843), .B(n99), .Q(n97) );
  NAND21 U492 ( .A(n823), .B(n192), .Q(n21) );
  AOI211 U493 ( .A(n822), .B(n857), .C(n856), .Q(n177) );
  AOI211 U494 ( .A(n822), .B(n167), .C(n168), .Q(n166) );
  XNR22 U495 ( .A(n21), .B(n193), .Q(SUM[14]) );
  INV2 U496 ( .A(n100), .Q(n850) );
  AOI211 U497 ( .A(n822), .B(n158), .C(n159), .Q(n157) );
  NAND20 U498 ( .A(n863), .B(n131), .Q(n14) );
  INV1 U500 ( .A(n131), .Q(n862) );
  AOI211 U501 ( .A(n840), .B(n90), .C(n91), .Q(n89) );
  OAI211 U502 ( .A(n176), .B(n802), .C(n177), .Q(n175) );
  NAND21 U503 ( .A(n841), .B(n145), .Q(n16) );
  NAND21 U504 ( .A(A[19]), .B(B[19]), .Q(n145) );
  OAI210 U505 ( .A(n92), .B(n850), .C(n95), .Q(n91) );
  XNR22 U506 ( .A(n9), .B(n87), .Q(SUM[26]) );
  NAND22 U507 ( .A(n825), .B(n167), .Q(n165) );
  INV3 U508 ( .A(n183), .Q(n825) );
  INV2 U509 ( .A(n244), .Q(n801) );
  XNR22 U510 ( .A(n7), .B(n69), .Q(SUM[28]) );
  BUF6 U512 ( .A(n141), .Q(n794) );
  BUF6 U513 ( .A(n123), .Q(n795) );
  NOR22 U514 ( .A(n81), .B(n115), .Q(n3) );
  NOR22 U515 ( .A(n149), .B(n183), .Q(n147) );
  NOR22 U516 ( .A(B[18]), .B(A[18]), .Q(n153) );
  INV0 U517 ( .A(n130), .Q(n863) );
  AOI211 U518 ( .A(n168), .B(n151), .C(n152), .Q(n150) );
  AOI212 U519 ( .A(n218), .B(n231), .C(n219), .Q(n217) );
  NAND20 U520 ( .A(n825), .B(n857), .Q(n176) );
  INV2 U521 ( .A(n156), .Q(n824) );
  INV0 U522 ( .A(n54), .Q(n812) );
  NAND21 U523 ( .A(n3), .B(n815), .Q(n59) );
  NAND22 U524 ( .A(n420), .B(n419), .Q(SUM[11]) );
  CLKIN3 U525 ( .A(n24), .Q(n847) );
  NAND20 U526 ( .A(n203), .B(n837), .Q(n194) );
  CLKIN0 U527 ( .A(n136), .Q(n839) );
  OAI210 U528 ( .A(n95), .B(n85), .C(n86), .Q(n84) );
  NAND21 U529 ( .A(n3), .B(n816), .Q(n70) );
  NAND22 U530 ( .A(n812), .B(n57), .Q(n6) );
  AOI210 U531 ( .A(n136), .B(n863), .C(n862), .Q(n127) );
  INV0 U532 ( .A(n405), .Q(n844) );
  NAND20 U533 ( .A(n135), .B(n863), .Q(n126) );
  NAND20 U534 ( .A(n815), .B(n45), .Q(n43) );
  INV0 U535 ( .A(n144), .Q(n841) );
  NAND20 U536 ( .A(n831), .B(n242), .Q(n28) );
  NOR20 U537 ( .A(n780), .B(n250), .Q(n245) );
  NAND20 U538 ( .A(n826), .B(n68), .Q(n7) );
  NAND20 U539 ( .A(n821), .B(n95), .Q(n10) );
  NAND21 U540 ( .A(n843), .B(n90), .Q(n88) );
  NAND20 U541 ( .A(n820), .B(n86), .Q(n9) );
  INV0 U542 ( .A(n105), .Q(n851) );
  AOI210 U543 ( .A(n62), .B(n45), .C(n46), .Q(n44) );
  INV0 U544 ( .A(n209), .Q(n845) );
  INV2 U545 ( .A(n67), .Q(n826) );
  INV0 U546 ( .A(n242), .Q(n829) );
  NAND20 U547 ( .A(A[24]), .B(B[24]), .Q(n106) );
  NOR20 U548 ( .A(B[4]), .B(A[4]), .Q(n254) );
  NAND20 U549 ( .A(A[26]), .B(B[26]), .Q(n86) );
  INV2 U550 ( .A(n74), .Q(n816) );
  NAND20 U551 ( .A(A[31]), .B(B[31]), .Q(n37) );
  NAND20 U552 ( .A(n3), .B(n810), .Q(n39) );
  NAND22 U553 ( .A(n707), .B(n844), .Q(n200) );
  NAND20 U554 ( .A(n802), .B(n847), .Q(n420) );
  NAND22 U555 ( .A(n200), .B(n22), .Q(n703) );
  INV3 U556 ( .A(n22), .Q(n836) );
  INV3 U557 ( .A(n411), .Q(n815) );
  NAND22 U558 ( .A(n843), .B(n855), .Q(n108) );
  INV3 U559 ( .A(n556), .Q(n819) );
  NAND22 U560 ( .A(n820), .B(n821), .Q(n556) );
  INV3 U561 ( .A(n43), .Q(n810) );
  INV3 U562 ( .A(n253), .Q(n800) );
  INV3 U563 ( .A(n265), .Q(n799) );
  NAND20 U564 ( .A(n828), .B(n781), .Q(n26) );
  AOI211 U565 ( .A(n801), .B(n230), .C(n779), .Q(n229) );
  NAND20 U566 ( .A(n827), .B(n221), .Q(n25) );
  AOI211 U567 ( .A(n801), .B(n223), .C(n224), .Q(n222) );
  XOR21 U568 ( .A(n30), .B(n800), .Q(SUM[5]) );
  NAND22 U569 ( .A(n859), .B(n251), .Q(n30) );
  INV2 U570 ( .A(n250), .Q(n859) );
  NAND20 U571 ( .A(n845), .B(n210), .Q(n23) );
  INV0 U572 ( .A(n191), .Q(n823) );
  NAND22 U573 ( .A(n846), .B(n124), .Q(n13) );
  INV3 U574 ( .A(n795), .Q(n846) );
  NAND22 U575 ( .A(n851), .B(n106), .Q(n11) );
  XNR21 U576 ( .A(n5), .B(n49), .Q(SUM[30]) );
  NAND22 U577 ( .A(n809), .B(n48), .Q(n5) );
  INV3 U578 ( .A(n47), .Q(n809) );
  XNR21 U579 ( .A(n29), .B(n249), .Q(SUM[6]) );
  XOR21 U580 ( .A(n256), .B(n31), .Q(SUM[4]) );
  NAND22 U581 ( .A(n807), .B(n255), .Q(n31) );
  INV3 U582 ( .A(n254), .Q(n807) );
  INV0 U583 ( .A(n168), .Q(n835) );
  INV1 U584 ( .A(n135), .Q(n842) );
  CLKIN3 U585 ( .A(n3), .Q(n818) );
  NAND22 U586 ( .A(n860), .B(n142), .Q(n15) );
  INV3 U587 ( .A(n794), .Q(n860) );
  NAND22 U588 ( .A(n853), .B(n163), .Q(n18) );
  NAND22 U589 ( .A(n833), .B(n174), .Q(n19) );
  INV3 U590 ( .A(n173), .Q(n833) );
  AOI211 U591 ( .A(n801), .B(n831), .C(n829), .Q(n238) );
  NOR21 U592 ( .A(n92), .B(n852), .Q(n90) );
  CLKIN3 U593 ( .A(n167), .Q(n834) );
  INV3 U594 ( .A(n75), .Q(n813) );
  AOI210 U595 ( .A(n2), .B(n810), .C(n811), .Q(n40) );
  INV3 U596 ( .A(n44), .Q(n811) );
  NAND20 U597 ( .A(n837), .B(n199), .Q(n22) );
  AOI211 U598 ( .A(n405), .B(n837), .C(n838), .Q(n195) );
  INV3 U599 ( .A(n181), .Q(n856) );
  NAND22 U601 ( .A(n826), .B(n816), .Q(n411) );
  NAND22 U602 ( .A(n858), .B(n154), .Q(n17) );
  NAND22 U603 ( .A(n700), .B(n157), .Q(n155) );
  INV3 U604 ( .A(n153), .Q(n858) );
  NAND22 U605 ( .A(n848), .B(n213), .Q(n24) );
  INV0 U606 ( .A(n212), .Q(n848) );
  INV3 U607 ( .A(n198), .Q(n837) );
  INV3 U608 ( .A(n112), .Q(n855) );
  INV3 U609 ( .A(n85), .Q(n820) );
  XOR21 U610 ( .A(n33), .B(n799), .Q(SUM[2]) );
  NAND22 U611 ( .A(n805), .B(n263), .Q(n33) );
  INV3 U612 ( .A(n262), .Q(n805) );
  XOR21 U613 ( .A(n269), .B(n34), .Q(SUM[1]) );
  NAND22 U614 ( .A(n804), .B(n267), .Q(n34) );
  INV3 U615 ( .A(n266), .Q(n804) );
  XNR21 U616 ( .A(n32), .B(n261), .Q(SUM[3]) );
  NAND22 U617 ( .A(n806), .B(n260), .Q(n32) );
  INV3 U618 ( .A(n259), .Q(n806) );
  AOI211 U619 ( .A(n265), .B(n257), .C(n258), .Q(n256) );
  NOR21 U620 ( .A(n259), .B(n262), .Q(n257) );
  XNR21 U621 ( .A(n4), .B(n38), .Q(SUM[31]) );
  NAND22 U622 ( .A(n808), .B(n37), .Q(n4) );
  NOR20 U624 ( .A(B[30]), .B(A[30]), .Q(n47) );
  NOR21 U625 ( .A(B[19]), .B(A[19]), .Q(n144) );
  NAND21 U626 ( .A(A[25]), .B(B[25]), .Q(n95) );
  NOR20 U627 ( .A(B[28]), .B(A[28]), .Q(n67) );
  NAND20 U628 ( .A(A[29]), .B(B[29]), .Q(n57) );
  NAND20 U629 ( .A(A[28]), .B(B[28]), .Q(n68) );
  NOR20 U630 ( .A(B[27]), .B(A[27]), .Q(n74) );
  NAND20 U631 ( .A(A[30]), .B(B[30]), .Q(n48) );
  INV3 U632 ( .A(n36), .Q(n808) );
  NOR20 U633 ( .A(B[31]), .B(A[31]), .Q(n36) );
  NAND20 U634 ( .A(A[4]), .B(B[4]), .Q(n255) );
  INV3 U635 ( .A(n35), .Q(SUM[0]) );
  NAND22 U636 ( .A(n798), .B(n269), .Q(n35) );
  INV3 U637 ( .A(n268), .Q(n798) );
  NOR20 U638 ( .A(B[0]), .B(A[0]), .Q(n268) );
  NOR20 U639 ( .A(B[3]), .B(A[3]), .Q(n259) );
  NOR20 U640 ( .A(B[2]), .B(A[2]), .Q(n262) );
  NAND20 U641 ( .A(A[0]), .B(B[0]), .Q(n269) );
  NAND20 U642 ( .A(A[2]), .B(B[2]), .Q(n263) );
  NOR20 U643 ( .A(B[1]), .B(A[1]), .Q(n266) );
  NAND20 U644 ( .A(A[1]), .B(B[1]), .Q(n267) );
  NAND20 U645 ( .A(A[3]), .B(B[3]), .Q(n260) );
  NOR21 U646 ( .A(B[5]), .B(A[5]), .Q(n250) );
  NAND22 U647 ( .A(A[12]), .B(B[12]), .Q(n210) );
  NOR23 U648 ( .A(B[14]), .B(A[14]), .Q(n191) );
  NAND20 U649 ( .A(n24), .B(n777), .Q(n419) );
  NOR21 U650 ( .A(B[21]), .B(A[21]), .Q(n130) );
endmodule


module adder_4 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_4_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n194,
         n195, n196, n197, n198, n203, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n420, n421, n427,
         n434, n435, n436, n440, n441, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  AOI212 U57 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  OAI212 U59 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U65 ( .A(n82), .B(n522), .C(n83), .Q(n81) );
  OAI212 U85 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  OAI212 U91 ( .A(n102), .B(n522), .C(n103), .Q(n101) );
  OAI212 U101 ( .A(n549), .B(n522), .C(n550), .Q(n108) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  AOI212 U107 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n522), .C(n159), .Q(n157) );
  OAI212 U175 ( .A(n585), .B(n522), .C(n583), .Q(n164) );
  OAI212 U183 ( .A(n177), .B(n173), .C(n174), .Q(n172) );
  OAI212 U197 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  AOI212 U249 ( .A(n221), .B(n240), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n527), .C(n227), .Q(n225) );
  OAI212 U275 ( .A(n245), .B(n241), .C(n242), .Q(n240) );
  OAI212 U281 ( .A(n518), .B(n527), .C(n245), .Q(n243) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  AOI212 U321 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U329 ( .A(n274), .B(n525), .C(n275), .Q(n273) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U423 ( .A(n252), .B(n256), .C(n253), .Q(n251) );
  OAI212 U464 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  AOI212 U412 ( .A(n526), .B(n258), .C(n427), .Q(n257) );
  OAI212 U401 ( .A(n120), .B(n522), .C(n121), .Q(n119) );
  OAI212 U405 ( .A(n129), .B(n522), .C(n130), .Q(n128) );
  OAI212 U525 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  OAI212 U413 ( .A(n64), .B(n522), .C(n65), .Q(n63) );
  OAI211 U349 ( .A(n73), .B(n522), .C(n74), .Q(n72) );
  OAI212 U350 ( .A(n188), .B(n527), .C(n189), .Q(n187) );
  NAND22 U351 ( .A(n261), .B(n571), .Q(n33) );
  INV0 U352 ( .A(n266), .Q(n591) );
  AOI212 U353 ( .A(n183), .B(n436), .C(n184), .Q(n182) );
  INV2 U354 ( .A(n436), .Q(n558) );
  INV3 U355 ( .A(n220), .Q(n562) );
  NOR23 U356 ( .A(n223), .B(n230), .Q(n221) );
  XOR22 U357 ( .A(n257), .B(n32), .Q(SUM[6]) );
  NAND21 U358 ( .A(n17), .B(n139), .Q(n420) );
  NAND23 U359 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NOR24 U360 ( .A(A[7]), .B(B[7]), .Q(n252) );
  NOR24 U361 ( .A(n252), .B(n255), .Q(n250) );
  NAND22 U362 ( .A(A[14]), .B(B[14]), .Q(n195) );
  NOR24 U363 ( .A(B[21]), .B(A[21]), .Q(n137) );
  INV2 U364 ( .A(n152), .Q(n577) );
  XNR22 U365 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NOR22 U366 ( .A(B[20]), .B(A[20]), .Q(n144) );
  NOR22 U367 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NAND23 U368 ( .A(n171), .B(n153), .Q(n151) );
  NOR23 U369 ( .A(n173), .B(n176), .Q(n171) );
  BUF15 U370 ( .A(n112), .Q(n506) );
  BUF2 U371 ( .A(n244), .Q(n518) );
  NAND22 U372 ( .A(A[10]), .B(B[10]), .Q(n231) );
  NOR21 U373 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR22 U374 ( .A(n155), .B(n162), .Q(n153) );
  NOR21 U375 ( .A(n70), .B(n6), .Q(n66) );
  NOR22 U376 ( .A(n137), .B(n144), .Q(n135) );
  NAND23 U377 ( .A(A[3]), .B(B[3]), .Q(n272) );
  INV3 U378 ( .A(n212), .Q(n573) );
  NAND23 U379 ( .A(n221), .B(n239), .Q(n219) );
  INV3 U380 ( .A(n219), .Q(n564) );
  NOR22 U381 ( .A(B[28]), .B(A[28]), .Q(n70) );
  NOR22 U382 ( .A(B[22]), .B(A[22]), .Q(n126) );
  NAND26 U383 ( .A(n511), .B(n512), .Q(SUM[19]) );
  NAND24 U384 ( .A(n509), .B(n510), .Q(n512) );
  INV3 U385 ( .A(n19), .Q(n509) );
  NAND24 U386 ( .A(n420), .B(n421), .Q(SUM[21]) );
  NAND22 U387 ( .A(n554), .B(n529), .Q(n421) );
  XOR21 U388 ( .A(n30), .B(n527), .Q(SUM[8]) );
  INV3 U389 ( .A(n23), .Q(n514) );
  NOR23 U390 ( .A(B[19]), .B(A[19]), .Q(n155) );
  BUF8 U391 ( .A(n111), .Q(n521) );
  OAI211 U392 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NAND21 U393 ( .A(n548), .B(n118), .Q(n15) );
  AOI210 U394 ( .A(n562), .B(n520), .C(n436), .Q(n198) );
  BUF2 U395 ( .A(n266), .Q(n507) );
  INV1 U396 ( .A(n562), .Q(n508) );
  NAND22 U397 ( .A(B[13]), .B(A[13]), .Q(n206) );
  NAND23 U398 ( .A(n203), .B(n183), .Q(n181) );
  NOR24 U399 ( .A(n185), .B(n194), .Q(n183) );
  NOR23 U400 ( .A(B[10]), .B(A[10]), .Q(n230) );
  NAND24 U402 ( .A(n514), .B(n515), .Q(n517) );
  INV3 U403 ( .A(n187), .Q(n515) );
  CLKIN4 U404 ( .A(n139), .Q(n529) );
  NOR23 U406 ( .A(B[8]), .B(A[8]), .Q(n244) );
  AOI212 U407 ( .A(n506), .B(n97), .C(n98), .Q(n92) );
  AOI212 U408 ( .A(n506), .B(n84), .C(n85), .Q(n83) );
  CLKIN2 U409 ( .A(n506), .Q(n550) );
  BUF6 U410 ( .A(n203), .Q(n520) );
  OAI212 U411 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  NOR22 U414 ( .A(n113), .B(n151), .Q(n111) );
  INV1 U415 ( .A(n117), .Q(n548) );
  INV0 U416 ( .A(n99), .Q(n545) );
  OAI212 U417 ( .A(n537), .B(n5), .C(n538), .Q(n56) );
  NAND22 U418 ( .A(n157), .B(n19), .Q(n511) );
  CLKIN6 U419 ( .A(n157), .Q(n510) );
  NAND22 U420 ( .A(n586), .B(n156), .Q(n19) );
  NAND24 U421 ( .A(A[8]), .B(B[8]), .Q(n245) );
  BUF15 U422 ( .A(n178), .Q(n522) );
  NAND21 U424 ( .A(n570), .B(n245), .Q(n30) );
  INV3 U425 ( .A(n566), .Q(n513) );
  CLKIN2 U426 ( .A(n240), .Q(n566) );
  OAI210 U427 ( .A(n260), .B(n266), .C(n261), .Q(n427) );
  NOR23 U428 ( .A(n265), .B(n260), .Q(n258) );
  INV0 U429 ( .A(n265), .Q(n590) );
  OAI212 U430 ( .A(n195), .B(n185), .C(n186), .Q(n184) );
  OAI211 U431 ( .A(n194), .B(n558), .C(n195), .Q(n191) );
  NAND28 U432 ( .A(n516), .B(n517), .Q(SUM[15]) );
  NAND22 U433 ( .A(A[18]), .B(B[18]), .Q(n163) );
  NOR22 U434 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NAND21 U435 ( .A(A[21]), .B(B[21]), .Q(n138) );
  CLKIN3 U436 ( .A(n230), .Q(n563) );
  NAND22 U437 ( .A(A[5]), .B(B[5]), .Q(n261) );
  NOR24 U438 ( .A(B[5]), .B(A[5]), .Q(n260) );
  INV1 U439 ( .A(n162), .Q(n575) );
  NAND22 U440 ( .A(n258), .B(n250), .Q(n248) );
  XOR21 U441 ( .A(n33), .B(n262), .Q(SUM[5]) );
  OAI212 U442 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  NOR22 U443 ( .A(n99), .B(n106), .Q(n97) );
  NOR24 U444 ( .A(B[13]), .B(A[13]), .Q(n205) );
  NAND22 U445 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NAND22 U446 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U447 ( .A(A[17]), .B(B[17]), .Q(n174) );
  AOI212 U448 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  NAND22 U449 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND22 U450 ( .A(n187), .B(n23), .Q(n516) );
  OAI212 U451 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  AOI211 U452 ( .A(n506), .B(n541), .C(n542), .Q(n74) );
  CLKIN4 U453 ( .A(n101), .Q(n528) );
  NOR22 U454 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NAND21 U455 ( .A(A[22]), .B(B[22]), .Q(n127) );
  NOR22 U456 ( .A(n181), .B(n219), .Q(n179) );
  OAI210 U457 ( .A(n42), .B(n522), .C(n43), .Q(n41) );
  NAND21 U458 ( .A(n580), .B(n253), .Q(n31) );
  NAND22 U459 ( .A(n175), .B(n21), .Q(n434) );
  NAND21 U460 ( .A(A[15]), .B(B[15]), .Q(n186) );
  NOR23 U461 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NOR23 U462 ( .A(B[12]), .B(A[12]), .Q(n212) );
  NAND22 U463 ( .A(n567), .B(n242), .Q(n29) );
  NAND22 U465 ( .A(B[9]), .B(A[9]), .Q(n242) );
  OAI211 U466 ( .A(n126), .B(n555), .C(n127), .Q(n123) );
  NOR24 U467 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NAND22 U468 ( .A(A[12]), .B(B[12]), .Q(n213) );
  OAI212 U469 ( .A(n197), .B(n527), .C(n198), .Q(n196) );
  NOR23 U470 ( .A(n79), .B(n519), .Q(n77) );
  NAND21 U471 ( .A(A[26]), .B(B[26]), .Q(n89) );
  NOR23 U472 ( .A(B[6]), .B(A[6]), .Q(n255) );
  XNR22 U473 ( .A(n8), .B(n52), .Q(SUM[30]) );
  CLKIN6 U474 ( .A(n175), .Q(n530) );
  NOR22 U475 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV8 U476 ( .A(n247), .Q(n527) );
  AOI211 U477 ( .A(n506), .B(n55), .C(n56), .Q(n54) );
  AOI211 U478 ( .A(n506), .B(n66), .C(n67), .Q(n65) );
  AOI212 U479 ( .A(n506), .B(n552), .C(n553), .Q(n103) );
  XNR21 U480 ( .A(n34), .B(n526), .Q(SUM[4]) );
  OAI212 U481 ( .A(n91), .B(n522), .C(n92), .Q(n90) );
  XNR22 U482 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U483 ( .A(n9), .B(n63), .Q(SUM[29]) );
  INV3 U484 ( .A(n255), .Q(n569) );
  INV4 U485 ( .A(n268), .Q(n526) );
  OAI212 U486 ( .A(n219), .B(n527), .C(n508), .Q(n214) );
  NOR21 U487 ( .A(B[24]), .B(A[24]), .Q(n106) );
  OAI211 U488 ( .A(n53), .B(n522), .C(n54), .Q(n52) );
  NAND21 U489 ( .A(n521), .B(n55), .Q(n53) );
  XNR22 U490 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI212 U491 ( .A(n151), .B(n522), .C(n152), .Q(n146) );
  NOR23 U492 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NOR24 U493 ( .A(B[11]), .B(A[11]), .Q(n223) );
  NAND21 U494 ( .A(B[11]), .B(A[11]), .Q(n224) );
  NAND22 U495 ( .A(n564), .B(n190), .Q(n188) );
  NOR22 U496 ( .A(n194), .B(n560), .Q(n190) );
  NOR20 U497 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR23 U498 ( .A(n205), .B(n212), .Q(n203) );
  OAI212 U499 ( .A(n260), .B(n266), .C(n261), .Q(n259) );
  NAND21 U500 ( .A(B[7]), .B(A[7]), .Q(n253) );
  INV0 U501 ( .A(n252), .Q(n580) );
  OAI212 U502 ( .A(n257), .B(n255), .C(n256), .Q(n254) );
  NOR23 U503 ( .A(n241), .B(n244), .Q(n239) );
  XNR22 U504 ( .A(n11), .B(n81), .Q(SUM[27]) );
  OAI212 U505 ( .A(n140), .B(n522), .C(n141), .Q(n139) );
  XNR22 U506 ( .A(n18), .B(n146), .Q(SUM[20]) );
  INV0 U507 ( .A(n205), .Q(n559) );
  XNR22 U508 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XNR22 U509 ( .A(n16), .B(n128), .Q(SUM[22]) );
  NAND24 U510 ( .A(n434), .B(n435), .Q(SUM[17]) );
  NAND22 U511 ( .A(n552), .B(n107), .Q(n14) );
  NAND21 U512 ( .A(A[24]), .B(B[24]), .Q(n107) );
  INV2 U513 ( .A(n5), .Q(n542) );
  OAI210 U514 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  NOR20 U515 ( .A(B[2]), .B(A[2]), .Q(n274) );
  XNR22 U516 ( .A(n27), .B(n225), .Q(SUM[11]) );
  AOI211 U517 ( .A(n526), .B(n590), .C(n591), .Q(n262) );
  XNR22 U518 ( .A(n26), .B(n214), .Q(SUM[12]) );
  XNR22 U519 ( .A(n20), .B(n164), .Q(SUM[18]) );
  NOR23 U520 ( .A(n117), .B(n126), .Q(n115) );
  NOR22 U521 ( .A(B[23]), .B(A[23]), .Q(n117) );
  CLKIN3 U522 ( .A(n163), .Q(n578) );
  NAND20 U523 ( .A(n575), .B(n163), .Q(n20) );
  OAI212 U524 ( .A(n208), .B(n527), .C(n209), .Q(n207) );
  OAI212 U526 ( .A(n176), .B(n522), .C(n177), .Q(n175) );
  OAI212 U527 ( .A(n568), .B(n527), .C(n566), .Q(n232) );
  INV2 U528 ( .A(n106), .Q(n552) );
  NAND23 U529 ( .A(n97), .B(n77), .Q(n6) );
  CLKIN3 U530 ( .A(n97), .Q(n546) );
  INV0 U531 ( .A(n173), .Q(n589) );
  NAND22 U532 ( .A(n521), .B(n541), .Q(n73) );
  XNR22 U533 ( .A(n243), .B(n29), .Q(SUM[9]) );
  XNR22 U534 ( .A(n24), .B(n196), .Q(SUM[14]) );
  XNR22 U535 ( .A(n25), .B(n207), .Q(SUM[13]) );
  NAND22 U536 ( .A(n521), .B(n552), .Q(n102) );
  NAND24 U537 ( .A(n440), .B(n441), .Q(SUM[25]) );
  NAND22 U538 ( .A(n576), .B(n135), .Q(n129) );
  NAND22 U539 ( .A(n576), .B(n122), .Q(n120) );
  NAND21 U540 ( .A(n576), .B(n582), .Q(n140) );
  INV2 U541 ( .A(n151), .Q(n576) );
  OAI212 U542 ( .A(n213), .B(n205), .C(n206), .Q(n436) );
  XNR22 U543 ( .A(n15), .B(n119), .Q(SUM[23]) );
  INV1 U544 ( .A(n185), .Q(n572) );
  AOI211 U545 ( .A(n562), .B(n190), .C(n191), .Q(n189) );
  XNR22 U546 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XOR21 U547 ( .A(n22), .B(n522), .Q(SUM[16]) );
  NAND21 U548 ( .A(n584), .B(n177), .Q(n22) );
  NAND21 U549 ( .A(n590), .B(n507), .Q(n34) );
  NAND21 U550 ( .A(n564), .B(n520), .Q(n197) );
  NAND22 U551 ( .A(n564), .B(n573), .Q(n208) );
  NAND21 U552 ( .A(n572), .B(n186), .Q(n23) );
  NAND22 U553 ( .A(n521), .B(n66), .Q(n64) );
  BUF6 U554 ( .A(n88), .Q(n519) );
  CLKIN3 U555 ( .A(n98), .Q(n547) );
  OAI212 U556 ( .A(n519), .B(n547), .C(n89), .Q(n85) );
  NOR21 U557 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NOR20 U558 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND21 U559 ( .A(n521), .B(n97), .Q(n91) );
  INV0 U560 ( .A(n176), .Q(n584) );
  CLKIN0 U561 ( .A(n171), .Q(n585) );
  CLKIN0 U562 ( .A(n172), .Q(n583) );
  NAND20 U563 ( .A(n551), .B(n127), .Q(n16) );
  CLKIN0 U564 ( .A(n135), .Q(n557) );
  NOR21 U565 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NAND20 U566 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV2 U567 ( .A(n21), .Q(n588) );
  NAND20 U568 ( .A(n171), .B(n575), .Q(n158) );
  NOR20 U569 ( .A(n46), .B(n6), .Q(n44) );
  NAND20 U570 ( .A(n239), .B(n563), .Q(n226) );
  CLKIN3 U571 ( .A(n59), .Q(n537) );
  CLKIN0 U572 ( .A(n239), .Q(n568) );
  AOI212 U573 ( .A(n250), .B(n259), .C(n251), .Q(n249) );
  INV0 U574 ( .A(n155), .Q(n586) );
  INV0 U575 ( .A(n126), .Q(n551) );
  NAND20 U576 ( .A(n563), .B(n231), .Q(n28) );
  CLKIN3 U577 ( .A(n521), .Q(n549) );
  INV0 U578 ( .A(n223), .Q(n579) );
  INV0 U579 ( .A(n194), .Q(n587) );
  CLKIN0 U580 ( .A(n144), .Q(n582) );
  INV0 U581 ( .A(n260), .Q(n571) );
  AOI210 U582 ( .A(n60), .B(n535), .C(n534), .Q(n47) );
  NAND20 U583 ( .A(n59), .B(n535), .Q(n46) );
  NAND20 U584 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U585 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U586 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U587 ( .A(A[27]), .B(B[27]), .Q(n80) );
  NAND20 U588 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NOR20 U589 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NOR21 U590 ( .A(n537), .B(n6), .Q(n55) );
  NAND20 U591 ( .A(n521), .B(n44), .Q(n42) );
  INV3 U592 ( .A(n6), .Q(n541) );
  INV3 U593 ( .A(n60), .Q(n538) );
  NAND22 U594 ( .A(n544), .B(n528), .Q(n441) );
  INV3 U595 ( .A(n13), .Q(n544) );
  AOI210 U596 ( .A(n577), .B(n135), .C(n136), .Q(n130) );
  INV3 U597 ( .A(n17), .Q(n554) );
  NAND22 U598 ( .A(n135), .B(n115), .Q(n113) );
  NAND22 U599 ( .A(n588), .B(n530), .Q(n435) );
  NAND22 U600 ( .A(n521), .B(n84), .Q(n82) );
  INV3 U601 ( .A(n277), .Q(n525) );
  NAND20 U602 ( .A(n569), .B(n256), .Q(n32) );
  INV3 U603 ( .A(n518), .Q(n570) );
  NAND22 U604 ( .A(n559), .B(n206), .Q(n25) );
  NAND20 U605 ( .A(n587), .B(n195), .Q(n24) );
  NAND20 U606 ( .A(n573), .B(n213), .Q(n26) );
  NAND22 U607 ( .A(n539), .B(n71), .Q(n10) );
  INV3 U608 ( .A(n70), .Q(n539) );
  NAND22 U609 ( .A(n536), .B(n62), .Q(n9) );
  INV3 U610 ( .A(n61), .Q(n536) );
  NAND22 U611 ( .A(n535), .B(n51), .Q(n8) );
  XNR21 U612 ( .A(n35), .B(n273), .Q(SUM[3]) );
  NAND22 U613 ( .A(n565), .B(n272), .Q(n35) );
  INV3 U614 ( .A(n271), .Q(n565) );
  NAND22 U615 ( .A(n543), .B(n89), .Q(n12) );
  INV3 U616 ( .A(n519), .Q(n543) );
  XOR21 U617 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND22 U618 ( .A(n531), .B(n279), .Q(n37) );
  INV3 U619 ( .A(n278), .Q(n531) );
  NOR21 U620 ( .A(n271), .B(n274), .Q(n269) );
  INV3 U621 ( .A(n520), .Q(n560) );
  AOI211 U622 ( .A(n577), .B(n582), .C(n581), .Q(n141) );
  INV3 U623 ( .A(n145), .Q(n581) );
  INV3 U624 ( .A(n51), .Q(n534) );
  INV3 U625 ( .A(n231), .Q(n561) );
  NAND22 U626 ( .A(n582), .B(n145), .Q(n18) );
  NAND22 U627 ( .A(n540), .B(n80), .Q(n11) );
  INV3 U628 ( .A(n79), .Q(n540) );
  NOR21 U629 ( .A(n61), .B(n70), .Q(n59) );
  INV0 U630 ( .A(n241), .Q(n567) );
  NAND20 U631 ( .A(n579), .B(n224), .Q(n27) );
  INV3 U632 ( .A(n107), .Q(n553) );
  NOR21 U633 ( .A(n519), .B(n546), .Q(n84) );
  AOI210 U634 ( .A(n172), .B(n575), .C(n578), .Q(n159) );
  AOI210 U635 ( .A(n577), .B(n122), .C(n123), .Q(n121) );
  CLKIN0 U636 ( .A(n136), .Q(n555) );
  NAND20 U637 ( .A(n589), .B(n174), .Q(n21) );
  AOI211 U638 ( .A(n562), .B(n573), .C(n574), .Q(n209) );
  INV0 U639 ( .A(n213), .Q(n574) );
  NAND20 U640 ( .A(n545), .B(n100), .Q(n13) );
  NAND20 U641 ( .A(n556), .B(n138), .Q(n17) );
  INV3 U642 ( .A(n137), .Q(n556) );
  NOR21 U643 ( .A(n126), .B(n557), .Q(n122) );
  XOR21 U644 ( .A(n36), .B(n525), .Q(SUM[2]) );
  NAND22 U645 ( .A(n532), .B(n275), .Q(n36) );
  INV3 U646 ( .A(n274), .Q(n532) );
  XNR21 U647 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U648 ( .A(n533), .B(n40), .Q(n7) );
  NAND21 U649 ( .A(A[19]), .B(B[19]), .Q(n156) );
  INV3 U650 ( .A(n50), .Q(n535) );
  NOR20 U651 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U652 ( .A(n39), .Q(n533) );
  INV3 U653 ( .A(n38), .Q(SUM[0]) );
  NAND22 U654 ( .A(n524), .B(n281), .Q(n38) );
  INV3 U655 ( .A(n280), .Q(n524) );
  NOR20 U656 ( .A(B[0]), .B(A[0]), .Q(n280) );
  NAND20 U657 ( .A(A[2]), .B(B[2]), .Q(n275) );
  NAND20 U658 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND20 U659 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NOR20 U660 ( .A(B[1]), .B(A[1]), .Q(n278) );
  NAND22 U661 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NAND22 U662 ( .A(n13), .B(n101), .Q(n440) );
  AOI210 U663 ( .A(n513), .B(n563), .C(n561), .Q(n227) );
  AOI210 U664 ( .A(n506), .B(n44), .C(n45), .Q(n43) );
endmodule


module adder_3 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_3_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n43, n44, n47, n48,
         n49, n50, n51, n52, n55, n56, n57, n58, n59, n60, n63, n64, n65, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n82, n83, n84,
         n85, n86, n87, n92, n93, n94, n95, n96, n99, n100, n101, n102, n103,
         n108, n109, n110, n111, n112, n113, n114, n117, n118, n119, n122,
         n123, n128, n129, n130, n131, n132, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n150, n151,
         n152, n153, n154, n155, n160, n161, n162, n163, n164, n167, n168,
         n169, n170, n171, n176, n177, n178, n179, n180, n181, n182, n185,
         n186, n187, n190, n191, n196, n197, n198, n199, n200, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n215, n216,
         n217, n218, n223, n224, n225, n228, n229, n231, n232, n233, n234,
         n235, n236, n237, n238, n240, n241, n242, n245, n246, n247, n250,
         n251, n253, n254, n255, n256, n257, n258, n259, n260, n262, n263,
         n264, n265, n266, n403, n404, n407, n408, n412, n418, n419, n422,
         n495, n499, n501, n506, n507, n582, n583, n594, n595, n598, n601,
         n602, n603, n760, n762, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943;

  OAI212 U48 ( .A(n68), .B(n103), .C(n69), .Q(n2) );
  AOI212 U100 ( .A(n123), .B(n108), .C(n109), .Q(n103) );
  OAI212 U118 ( .A(n911), .B(n864), .C(n910), .Q(n119) );
  OAI212 U126 ( .A(n132), .B(n412), .C(n129), .Q(n123) );
  AOI212 U138 ( .A(n202), .B(n134), .C(n135), .Q(n1) );
  OAI212 U231 ( .A(n203), .B(n231), .C(n204), .Q(n202) );
  OAI212 U287 ( .A(n241), .B(n253), .C(n242), .Q(n240) );
  OAI212 U308 ( .A(n260), .B(n256), .C(n257), .Q(n255) );
  OAI212 U314 ( .A(n259), .B(n934), .C(n260), .Q(n258) );
  OAI212 U321 ( .A(n266), .B(n263), .C(n264), .Q(n262) );
  OAI212 U414 ( .A(n118), .B(n603), .C(n111), .Q(n109) );
  OAI212 U443 ( .A(n422), .B(n864), .C(n132), .Q(n130) );
  OAI212 U458 ( .A(n113), .B(n864), .C(n114), .Q(n112) );
  OAI212 U619 ( .A(n95), .B(n864), .C(n96), .Q(n94) );
  OAI212 U409 ( .A(n75), .B(n864), .C(n76), .Q(n74) );
  OAI212 U450 ( .A(n84), .B(n864), .C(n85), .Q(n83) );
  OAI212 U339 ( .A(n59), .B(n864), .C(n60), .Q(n58) );
  OAI212 U353 ( .A(n872), .B(n864), .C(n869), .Q(n65) );
  OAI212 U412 ( .A(n922), .B(n918), .C(n923), .Q(n187) );
  OAI212 U423 ( .A(n181), .B(n918), .C(n182), .Q(n180) );
  OAI212 U397 ( .A(n936), .B(n237), .C(n238), .Q(n236) );
  AOI212 U435 ( .A(n205), .B(n501), .C(n206), .Q(n204) );
  OAI212 U463 ( .A(n168), .B(n160), .C(n161), .Q(n155) );
  OAI212 U386 ( .A(n39), .B(n864), .C(n40), .Q(n38) );
  OAI212 U431 ( .A(n171), .B(n136), .C(n137), .Q(n135) );
  OAI212 U491 ( .A(n143), .B(n918), .C(n144), .Q(n142) );
  OAI212 U352 ( .A(n422), .B(n864), .C(n132), .Q(n760) );
  OAI212 U417 ( .A(n64), .B(n56), .C(n57), .Q(n55) );
  OAI212 U510 ( .A(n859), .B(n919), .C(n215), .Q(n211) );
  CLKIN3 U334 ( .A(n119), .Q(n898) );
  NAND24 U335 ( .A(n582), .B(n583), .Q(SUM[27]) );
  INV2 U336 ( .A(n2), .Q(n869) );
  INV6 U337 ( .A(n94), .Q(n883) );
  NOR22 U338 ( .A(n128), .B(n131), .Q(n122) );
  INV6 U340 ( .A(n102), .Q(n891) );
  NAND22 U341 ( .A(n101), .B(n11), .Q(n601) );
  NOR23 U342 ( .A(A[16]), .B(B[16]), .Q(n167) );
  CLKIN6 U343 ( .A(n130), .Q(n899) );
  NAND23 U344 ( .A(n86), .B(n70), .Q(n68) );
  NAND21 U345 ( .A(A[21]), .B(B[21]), .Q(n129) );
  NAND24 U346 ( .A(n854), .B(n855), .Q(SUM[19]) );
  NAND24 U347 ( .A(n852), .B(n853), .Q(n855) );
  NOR24 U348 ( .A(A[17]), .B(B[17]), .Q(n160) );
  XNR22 U349 ( .A(n17), .B(n151), .Q(SUM[18]) );
  NAND26 U350 ( .A(n850), .B(n851), .Q(SUM[13]) );
  NAND24 U351 ( .A(n848), .B(n849), .Q(n851) );
  XNR22 U354 ( .A(n19), .B(n169), .Q(SUM[16]) );
  NAND22 U355 ( .A(A[11]), .B(B[11]), .Q(n208) );
  NOR21 U356 ( .A(B[22]), .B(A[22]), .Q(n117) );
  CLKIN4 U357 ( .A(n101), .Q(n890) );
  OAI212 U358 ( .A(n102), .B(n864), .C(n103), .Q(n101) );
  NOR24 U359 ( .A(n110), .B(n857), .Q(n108) );
  BUF15 U360 ( .A(n167), .Q(n863) );
  NAND26 U361 ( .A(n601), .B(n602), .Q(SUM[24]) );
  AOI212 U362 ( .A(n904), .B(n145), .C(n146), .Q(n144) );
  NOR24 U363 ( .A(n92), .B(n99), .Q(n86) );
  NOR22 U364 ( .A(B[24]), .B(A[24]), .Q(n99) );
  NAND22 U365 ( .A(A[16]), .B(B[16]), .Q(n168) );
  NOR24 U366 ( .A(B[9]), .B(A[9]), .Q(n223) );
  NAND24 U367 ( .A(B[9]), .B(A[9]), .Q(n224) );
  NOR22 U368 ( .A(n136), .B(n170), .Q(n134) );
  INV3 U369 ( .A(n142), .Q(n853) );
  INV3 U370 ( .A(n112), .Q(n892) );
  NOR22 U371 ( .A(B[18]), .B(A[18]), .Q(n495) );
  NAND22 U372 ( .A(A[18]), .B(B[18]), .Q(n150) );
  INV3 U373 ( .A(n198), .Q(n848) );
  NOR22 U374 ( .A(n856), .B(n79), .Q(n70) );
  NOR21 U375 ( .A(B[26]), .B(A[26]), .Q(n79) );
  AOI211 U376 ( .A(n232), .B(n240), .C(n233), .Q(n231) );
  INV3 U377 ( .A(n74), .Q(n877) );
  NAND24 U378 ( .A(n893), .B(n898), .Q(n419) );
  INV3 U379 ( .A(n160), .Q(n928) );
  NAND26 U380 ( .A(n594), .B(n595), .Q(SUM[25]) );
  NAND24 U381 ( .A(n878), .B(n883), .Q(n595) );
  NAND26 U382 ( .A(n407), .B(n408), .Q(SUM[21]) );
  NAND24 U383 ( .A(n403), .B(n404), .Q(SUM[23]) );
  NAND23 U384 ( .A(n887), .B(n892), .Q(n404) );
  AOI211 U385 ( .A(n921), .B(n217), .C(n218), .Q(n216) );
  XOR21 U387 ( .A(n24), .B(n209), .Q(SUM[11]) );
  INV3 U388 ( .A(n207), .Q(n927) );
  INV3 U389 ( .A(n22), .Q(n849) );
  NAND22 U390 ( .A(n902), .B(n186), .Q(n21) );
  INV3 U391 ( .A(n904), .Q(n847) );
  NOR22 U392 ( .A(B[25]), .B(A[25]), .Q(n92) );
  NAND21 U393 ( .A(n122), .B(n894), .Q(n113) );
  INV1 U394 ( .A(n155), .Q(n901) );
  NOR22 U395 ( .A(n68), .B(n102), .Q(n3) );
  OAI211 U396 ( .A(n238), .B(n234), .C(n235), .Q(n233) );
  NAND26 U398 ( .A(n418), .B(n419), .Q(SUM[22]) );
  OAI212 U399 ( .A(n200), .B(n196), .C(n197), .Q(n191) );
  AOI211 U400 ( .A(n2), .B(n52), .C(n55), .Q(n51) );
  NAND22 U401 ( .A(A[19]), .B(B[19]), .Q(n141) );
  NAND21 U402 ( .A(n927), .B(n208), .Q(n24) );
  NOR22 U403 ( .A(B[10]), .B(A[10]), .Q(n212) );
  NOR22 U404 ( .A(n207), .B(n212), .Q(n205) );
  XOR22 U405 ( .A(n25), .B(n216), .Q(SUM[10]) );
  CLKIN0 U406 ( .A(n168), .Q(n900) );
  INV1 U407 ( .A(n185), .Q(n902) );
  NAND24 U408 ( .A(n190), .B(n176), .Q(n170) );
  NOR20 U410 ( .A(A[28]), .B(B[28]), .Q(n63) );
  NOR21 U411 ( .A(B[23]), .B(A[23]), .Q(n110) );
  NAND26 U413 ( .A(n875), .B(n881), .Q(n507) );
  NAND22 U415 ( .A(n198), .B(n22), .Q(n850) );
  NAND24 U416 ( .A(n862), .B(n200), .Q(n198) );
  NAND22 U418 ( .A(n931), .B(n197), .Q(n22) );
  NOR20 U419 ( .A(A[30]), .B(B[30]), .Q(n47) );
  OAI211 U420 ( .A(n113), .B(n864), .C(n114), .Q(n762) );
  NAND22 U421 ( .A(n16), .B(n142), .Q(n854) );
  INV2 U422 ( .A(n16), .Q(n852) );
  AOI212 U424 ( .A(n87), .B(n70), .C(n71), .Q(n69) );
  NAND22 U425 ( .A(n8), .B(n74), .Q(n582) );
  NAND22 U426 ( .A(n9), .B(n83), .Q(n506) );
  NAND28 U427 ( .A(n506), .B(n507), .Q(SUM[26]) );
  INV6 U428 ( .A(n103), .Q(n889) );
  NAND20 U429 ( .A(n909), .B(n129), .Q(n14) );
  NOR24 U430 ( .A(B[11]), .B(A[11]), .Q(n207) );
  NAND22 U432 ( .A(B[14]), .B(A[14]), .Q(n186) );
  NOR23 U433 ( .A(A[15]), .B(B[15]), .Q(n178) );
  NOR23 U434 ( .A(n196), .B(n199), .Q(n190) );
  OAI212 U436 ( .A(n100), .B(n92), .C(n93), .Q(n87) );
  NAND21 U437 ( .A(A[24]), .B(B[24]), .Q(n100) );
  NAND28 U438 ( .A(A[8]), .B(B[8]), .Q(n229) );
  NOR21 U439 ( .A(B[8]), .B(A[8]), .Q(n228) );
  NOR21 U440 ( .A(n223), .B(n228), .Q(n217) );
  OAI212 U441 ( .A(n229), .B(n223), .C(n224), .Q(n218) );
  INV2 U442 ( .A(n223), .Q(n916) );
  CLKIN12 U444 ( .A(n202), .Q(n918) );
  INV6 U445 ( .A(n918), .Q(n861) );
  AOI211 U446 ( .A(n889), .B(n77), .C(n78), .Q(n76) );
  NAND24 U447 ( .A(n870), .B(n877), .Q(n583) );
  OAI211 U448 ( .A(n79), .B(n882), .C(n82), .Q(n78) );
  AOI212 U449 ( .A(n155), .B(n138), .C(n139), .Q(n137) );
  OAI211 U451 ( .A(n163), .B(n918), .C(n164), .Q(n162) );
  INV3 U452 ( .A(n171), .Q(n904) );
  NAND24 U453 ( .A(n154), .B(n138), .Q(n136) );
  INV2 U454 ( .A(n154), .Q(n897) );
  NOR20 U455 ( .A(B[10]), .B(A[10]), .Q(n859) );
  NAND23 U456 ( .A(A[10]), .B(B[10]), .Q(n215) );
  NAND22 U457 ( .A(n119), .B(n13), .Q(n418) );
  INV0 U459 ( .A(n186), .Q(n905) );
  AOI211 U460 ( .A(n904), .B(n154), .C(n155), .Q(n153) );
  OAI211 U461 ( .A(n152), .B(n918), .C(n153), .Q(n151) );
  NOR21 U462 ( .A(B[23]), .B(A[23]), .Q(n603) );
  OAI211 U464 ( .A(n82), .B(n856), .C(n73), .Q(n71) );
  NOR23 U465 ( .A(B[19]), .B(A[19]), .Q(n140) );
  NOR23 U466 ( .A(n140), .B(n147), .Q(n138) );
  INV6 U467 ( .A(n170), .Q(n903) );
  NOR21 U468 ( .A(B[6]), .B(A[6]), .Q(n237) );
  XNR22 U469 ( .A(n6), .B(n58), .Q(SUM[29]) );
  CLKIN6 U470 ( .A(n83), .Q(n881) );
  NAND22 U471 ( .A(n94), .B(n10), .Q(n594) );
  NOR21 U472 ( .A(B[21]), .B(A[21]), .Q(n412) );
  OAI211 U473 ( .A(n50), .B(n864), .C(n51), .Q(n49) );
  CLKIN2 U474 ( .A(n140), .Q(n912) );
  OAI212 U475 ( .A(n229), .B(n223), .C(n224), .Q(n501) );
  XNR22 U476 ( .A(n21), .B(n187), .Q(SUM[14]) );
  NAND22 U477 ( .A(n929), .B(n179), .Q(n20) );
  NAND21 U478 ( .A(A[15]), .B(B[15]), .Q(n179) );
  NAND21 U479 ( .A(n891), .B(n86), .Q(n84) );
  NAND24 U480 ( .A(n885), .B(n890), .Q(n602) );
  NAND26 U481 ( .A(n899), .B(n908), .Q(n408) );
  NAND24 U482 ( .A(A[12]), .B(B[12]), .Q(n200) );
  NAND21 U483 ( .A(A[17]), .B(B[17]), .Q(n161) );
  XOR22 U484 ( .A(n15), .B(n864), .Q(SUM[20]) );
  NAND20 U485 ( .A(n886), .B(n100), .Q(n11) );
  CLKIN3 U486 ( .A(n87), .Q(n882) );
  AOI211 U487 ( .A(n889), .B(n86), .C(n87), .Q(n85) );
  OAI212 U488 ( .A(n186), .B(n178), .C(n179), .Q(n177) );
  NAND22 U489 ( .A(n3), .B(n52), .Q(n50) );
  NOR23 U490 ( .A(n178), .B(n185), .Q(n176) );
  NOR22 U492 ( .A(B[14]), .B(A[14]), .Q(n185) );
  XNR22 U493 ( .A(n20), .B(n180), .Q(SUM[15]) );
  NOR22 U494 ( .A(B[18]), .B(A[18]), .Q(n147) );
  BUF15 U495 ( .A(n1), .Q(n864) );
  XNR22 U496 ( .A(n18), .B(n162), .Q(SUM[17]) );
  XNR22 U497 ( .A(n7), .B(n65), .Q(SUM[28]) );
  INV1 U498 ( .A(n100), .Q(n884) );
  OAI211 U499 ( .A(n901), .B(n495), .C(n150), .Q(n146) );
  NAND21 U500 ( .A(n916), .B(n224), .Q(n26) );
  OAI212 U501 ( .A(n215), .B(n207), .C(n208), .Q(n206) );
  NAND22 U502 ( .A(A[20]), .B(B[20]), .Q(n132) );
  NOR24 U503 ( .A(A[13]), .B(B[13]), .Q(n196) );
  BUF6 U504 ( .A(n72), .Q(n856) );
  OAI211 U505 ( .A(n170), .B(n918), .C(n847), .Q(n169) );
  AOI212 U506 ( .A(n191), .B(n176), .C(n177), .Q(n171) );
  BUF6 U507 ( .A(n117), .Q(n857) );
  NOR24 U508 ( .A(n160), .B(n863), .Q(n154) );
  NAND24 U509 ( .A(A[13]), .B(B[13]), .Q(n197) );
  NOR20 U511 ( .A(B[10]), .B(A[10]), .Q(n858) );
  NAND24 U512 ( .A(n860), .B(n861), .Q(n862) );
  INV0 U513 ( .A(n199), .Q(n860) );
  NOR22 U514 ( .A(B[12]), .B(A[12]), .Q(n199) );
  CLKIN1 U515 ( .A(n86), .Q(n880) );
  NAND22 U516 ( .A(n145), .B(n903), .Q(n143) );
  NAND22 U517 ( .A(n860), .B(n200), .Q(n23) );
  INV0 U518 ( .A(n858), .Q(n924) );
  OAI210 U519 ( .A(n200), .B(n196), .C(n197), .Q(n499) );
  CLKIN2 U520 ( .A(n10), .Q(n878) );
  NAND22 U521 ( .A(n891), .B(n886), .Q(n95) );
  AOI211 U522 ( .A(n889), .B(n886), .C(n884), .Q(n96) );
  CLKIN0 U523 ( .A(n122), .Q(n911) );
  INV2 U524 ( .A(n13), .Q(n893) );
  CLKIN3 U525 ( .A(n9), .Q(n875) );
  INV0 U526 ( .A(n123), .Q(n910) );
  INV0 U527 ( .A(n196), .Q(n931) );
  CLKIN2 U528 ( .A(n499), .Q(n923) );
  CLKIN3 U529 ( .A(n218), .Q(n919) );
  CLKIN0 U530 ( .A(n190), .Q(n922) );
  NAND20 U531 ( .A(n896), .B(n168), .Q(n19) );
  NAND21 U532 ( .A(A[22]), .B(B[22]), .Q(n118) );
  NAND20 U533 ( .A(A[4]), .B(B[4]), .Q(n251) );
  NAND20 U534 ( .A(A[5]), .B(B[5]), .Q(n246) );
  NAND20 U535 ( .A(n903), .B(n154), .Q(n152) );
  NAND20 U536 ( .A(n903), .B(n896), .Q(n163) );
  NAND20 U537 ( .A(n912), .B(n141), .Q(n16) );
  INV0 U538 ( .A(n178), .Q(n929) );
  NAND20 U539 ( .A(n894), .B(n118), .Q(n13) );
  NOR20 U540 ( .A(B[27]), .B(A[27]), .Q(n72) );
  NOR20 U541 ( .A(B[20]), .B(A[20]), .Q(n131) );
  NOR20 U542 ( .A(B[21]), .B(A[21]), .Q(n128) );
  NAND20 U543 ( .A(n217), .B(n205), .Q(n203) );
  NOR20 U544 ( .A(B[20]), .B(A[20]), .Q(n422) );
  NAND20 U545 ( .A(A[26]), .B(B[26]), .Q(n82) );
  NAND20 U546 ( .A(A[25]), .B(B[25]), .Q(n93) );
  NAND20 U547 ( .A(A[27]), .B(B[27]), .Q(n73) );
  NAND20 U548 ( .A(A[23]), .B(B[23]), .Q(n111) );
  INV2 U549 ( .A(n237), .Q(n930) );
  NOR21 U550 ( .A(n56), .B(n63), .Q(n52) );
  NOR20 U551 ( .A(n234), .B(n237), .Q(n232) );
  NAND20 U552 ( .A(B[28]), .B(A[28]), .Q(n64) );
  NOR20 U553 ( .A(B[7]), .B(A[7]), .Q(n234) );
  NAND20 U554 ( .A(B[30]), .B(A[30]), .Q(n48) );
  NAND22 U555 ( .A(n762), .B(n12), .Q(n403) );
  INV3 U556 ( .A(n11), .Q(n885) );
  INV3 U557 ( .A(n8), .Q(n870) );
  NAND22 U558 ( .A(n190), .B(n902), .Q(n181) );
  INV3 U559 ( .A(n14), .Q(n908) );
  INV3 U560 ( .A(n12), .Q(n887) );
  NAND22 U561 ( .A(n891), .B(n77), .Q(n75) );
  NOR21 U562 ( .A(n79), .B(n880), .Q(n77) );
  NAND22 U563 ( .A(n913), .B(n132), .Q(n15) );
  INV3 U564 ( .A(n422), .Q(n913) );
  NAND22 U565 ( .A(n924), .B(n215), .Q(n25) );
  XOR21 U566 ( .A(n26), .B(n225), .Q(SUM[9]) );
  AOI211 U567 ( .A(n921), .B(n925), .C(n926), .Q(n225) );
  INV3 U568 ( .A(n229), .Q(n926) );
  XOR21 U569 ( .A(n23), .B(n918), .Q(SUM[12]) );
  XNR21 U570 ( .A(n27), .B(n921), .Q(SUM[8]) );
  NAND22 U571 ( .A(n925), .B(n229), .Q(n27) );
  NAND22 U572 ( .A(n928), .B(n161), .Q(n18) );
  NAND22 U573 ( .A(n915), .B(n150), .Q(n17) );
  INV3 U574 ( .A(n495), .Q(n915) );
  AOI210 U575 ( .A(n123), .B(n894), .C(n895), .Q(n114) );
  INV3 U576 ( .A(n118), .Q(n895) );
  AOI211 U577 ( .A(n921), .B(n210), .C(n211), .Q(n209) );
  NAND22 U578 ( .A(n122), .B(n108), .Q(n102) );
  NAND22 U579 ( .A(n879), .B(n93), .Q(n10) );
  INV3 U580 ( .A(n92), .Q(n879) );
  INV3 U581 ( .A(n412), .Q(n909) );
  NAND22 U582 ( .A(n111), .B(n888), .Q(n12) );
  INV3 U583 ( .A(n603), .Q(n888) );
  NOR21 U584 ( .A(n495), .B(n897), .Q(n145) );
  NAND22 U585 ( .A(n598), .B(n141), .Q(n139) );
  NAND22 U586 ( .A(n914), .B(n912), .Q(n598) );
  INV3 U587 ( .A(n150), .Q(n914) );
  NAND22 U588 ( .A(n876), .B(n82), .Q(n9) );
  INV3 U589 ( .A(n79), .Q(n876) );
  NAND22 U590 ( .A(n871), .B(n73), .Q(n8) );
  INV3 U591 ( .A(n856), .Q(n871) );
  AOI211 U592 ( .A(n904), .B(n896), .C(n900), .Q(n164) );
  AOI211 U593 ( .A(n499), .B(n902), .C(n905), .Q(n182) );
  NAND22 U594 ( .A(n760), .B(n14), .Q(n407) );
  INV3 U595 ( .A(n857), .Q(n894) );
  INV3 U596 ( .A(n863), .Q(n896) );
  INV3 U597 ( .A(n99), .Q(n886) );
  INV3 U598 ( .A(n228), .Q(n925) );
  NOR21 U599 ( .A(n858), .B(n917), .Q(n210) );
  INV3 U600 ( .A(n217), .Q(n917) );
  NAND22 U601 ( .A(n3), .B(n873), .Q(n59) );
  NAND20 U602 ( .A(n3), .B(n868), .Q(n39) );
  INV3 U603 ( .A(n231), .Q(n921) );
  INV3 U604 ( .A(n240), .Q(n936) );
  INV3 U605 ( .A(n262), .Q(n934) );
  INV3 U606 ( .A(n253), .Q(n935) );
  NAND22 U607 ( .A(n867), .B(n57), .Q(n6) );
  CLKIN3 U608 ( .A(n56), .Q(n867) );
  NAND22 U609 ( .A(n873), .B(n64), .Q(n7) );
  INV3 U610 ( .A(n3), .Q(n872) );
  XNR21 U611 ( .A(n5), .B(n49), .Q(SUM[30]) );
  NAND22 U612 ( .A(n906), .B(n48), .Q(n5) );
  XNR21 U613 ( .A(n28), .B(n236), .Q(SUM[7]) );
  NAND22 U614 ( .A(n920), .B(n235), .Q(n28) );
  INV3 U615 ( .A(n234), .Q(n920) );
  XOR21 U616 ( .A(n936), .B(n29), .Q(SUM[6]) );
  NAND22 U617 ( .A(n930), .B(n238), .Q(n29) );
  CLKIN3 U618 ( .A(n63), .Q(n873) );
  AOI211 U620 ( .A(n2), .B(n873), .C(n874), .Q(n60) );
  INV3 U621 ( .A(n64), .Q(n874) );
  AOI210 U622 ( .A(n2), .B(n868), .C(n866), .Q(n40) );
  CLKIN3 U623 ( .A(n44), .Q(n866) );
  AOI210 U624 ( .A(n55), .B(n906), .C(n907), .Q(n44) );
  INV3 U625 ( .A(n48), .Q(n907) );
  INV3 U626 ( .A(n43), .Q(n868) );
  NAND20 U627 ( .A(n52), .B(n906), .Q(n43) );
  XOR21 U628 ( .A(n30), .B(n247), .Q(SUM[5]) );
  NAND22 U629 ( .A(n943), .B(n246), .Q(n30) );
  AOI211 U630 ( .A(n935), .B(n941), .C(n940), .Q(n247) );
  XOR21 U631 ( .A(n33), .B(n934), .Q(SUM[2]) );
  NAND22 U632 ( .A(n938), .B(n260), .Q(n33) );
  INV3 U633 ( .A(n259), .Q(n938) );
  XOR21 U634 ( .A(n266), .B(n34), .Q(SUM[1]) );
  NAND22 U635 ( .A(n937), .B(n264), .Q(n34) );
  INV3 U636 ( .A(n263), .Q(n937) );
  NAND22 U637 ( .A(n941), .B(n943), .Q(n241) );
  AOI211 U638 ( .A(n943), .B(n940), .C(n942), .Q(n242) );
  INV3 U639 ( .A(n246), .Q(n942) );
  XNR21 U640 ( .A(n32), .B(n258), .Q(SUM[3]) );
  NAND22 U641 ( .A(n939), .B(n257), .Q(n32) );
  INV3 U642 ( .A(n256), .Q(n939) );
  AOI211 U643 ( .A(n262), .B(n254), .C(n255), .Q(n253) );
  NOR21 U644 ( .A(n256), .B(n259), .Q(n254) );
  XNR21 U645 ( .A(n31), .B(n935), .Q(SUM[4]) );
  NAND22 U646 ( .A(n941), .B(n251), .Q(n31) );
  INV3 U647 ( .A(n251), .Q(n940) );
  XNR21 U648 ( .A(n4), .B(n38), .Q(SUM[31]) );
  NAND22 U649 ( .A(n865), .B(n37), .Q(n4) );
  NAND20 U650 ( .A(B[31]), .B(A[31]), .Q(n37) );
  NAND20 U651 ( .A(B[29]), .B(A[29]), .Q(n57) );
  INV3 U652 ( .A(n47), .Q(n906) );
  INV3 U653 ( .A(n36), .Q(n865) );
  NAND20 U654 ( .A(A[6]), .B(B[6]), .Q(n238) );
  NAND20 U655 ( .A(A[7]), .B(B[7]), .Q(n235) );
  INV3 U656 ( .A(n245), .Q(n943) );
  NOR20 U657 ( .A(B[5]), .B(A[5]), .Q(n245) );
  INV3 U658 ( .A(n35), .Q(SUM[0]) );
  NAND22 U659 ( .A(n933), .B(n266), .Q(n35) );
  INV3 U660 ( .A(n265), .Q(n933) );
  NOR20 U661 ( .A(B[0]), .B(A[0]), .Q(n265) );
  INV3 U662 ( .A(n250), .Q(n941) );
  NOR20 U663 ( .A(B[4]), .B(A[4]), .Q(n250) );
  NOR20 U664 ( .A(B[3]), .B(A[3]), .Q(n256) );
  NOR20 U665 ( .A(B[2]), .B(A[2]), .Q(n259) );
  NAND20 U666 ( .A(A[0]), .B(B[0]), .Q(n266) );
  NAND20 U667 ( .A(A[2]), .B(B[2]), .Q(n260) );
  NOR20 U668 ( .A(B[1]), .B(A[1]), .Q(n263) );
  NAND20 U669 ( .A(A[1]), .B(B[1]), .Q(n264) );
  NAND20 U670 ( .A(A[3]), .B(B[3]), .Q(n257) );
  NOR21 U671 ( .A(A[31]), .B(B[31]), .Q(n36) );
  NOR21 U672 ( .A(A[29]), .B(B[29]), .Q(n56) );
endmodule


module adder_2 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_2_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module adder_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n88, n89, n90, n91, n92, n97, n98, n99, n100, n101, n102,
         n103, n106, n107, n108, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n126, n127, n128, n129, n130,
         n135, n136, n137, n138, n139, n140, n141, n144, n145, n146, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n230, n231, n232, n239, n240, n241, n242, n243, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n265, n266, n268, n269, n270, n271, n272,
         n273, n274, n275, n277, n278, n279, n280, n281, n418, n419, n424,
         n425, n430, n431, n436, n437, n438, n444, n448, n449, n450, n455,
         n456, n461, n462, n463, n470, n471, n472, n473, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645;

  OAI212 U77 ( .A(n91), .B(n566), .C(n92), .Q(n90) );
  OAI212 U105 ( .A(n113), .B(n152), .C(n114), .Q(n112) );
  OAI212 U115 ( .A(n120), .B(n566), .C(n121), .Q(n119) );
  OAI212 U127 ( .A(n129), .B(n566), .C(n130), .Q(n128) );
  OAI212 U141 ( .A(n140), .B(n566), .C(n141), .Q(n139) );
  OAI212 U151 ( .A(n151), .B(n566), .C(n463), .Q(n146) );
  AOI212 U157 ( .A(n172), .B(n153), .C(n154), .Q(n152) );
  OAI212 U165 ( .A(n158), .B(n566), .C(n159), .Q(n157) );
  OAI212 U183 ( .A(n173), .B(n177), .C(n174), .Q(n172) );
  OAI212 U189 ( .A(n176), .B(n566), .C(n177), .Q(n175) );
  AOI212 U195 ( .A(n247), .B(n179), .C(n180), .Q(n178) );
  OAI212 U219 ( .A(n197), .B(n584), .C(n198), .Q(n196) );
  AOI212 U249 ( .A(n240), .B(n221), .C(n222), .Q(n220) );
  OAI212 U251 ( .A(n231), .B(n223), .C(n224), .Q(n222) );
  OAI212 U257 ( .A(n226), .B(n584), .C(n227), .Q(n225) );
  OAI212 U267 ( .A(n581), .B(n584), .C(n578), .Q(n232) );
  OAI212 U288 ( .A(n248), .B(n268), .C(n249), .Q(n247) );
  AOI212 U290 ( .A(n259), .B(n250), .C(n251), .Q(n249) );
  AOI212 U321 ( .A(n277), .B(n269), .C(n270), .Q(n268) );
  OAI212 U336 ( .A(n281), .B(n278), .C(n279), .Q(n277) );
  OAI212 U391 ( .A(n107), .B(n99), .C(n100), .Q(n98) );
  AOI212 U433 ( .A(n136), .B(n115), .C(n116), .Q(n114) );
  OAI212 U512 ( .A(n145), .B(n137), .C(n138), .Q(n136) );
  XOR22 U489 ( .A(n22), .B(n566), .Q(SUM[16]) );
  OAI212 U500 ( .A(n127), .B(n117), .C(n118), .Q(n116) );
  AOI212 U354 ( .A(n588), .B(n589), .C(n590), .Q(n262) );
  NOR24 U379 ( .A(n205), .B(n212), .Q(n203) );
  OAI212 U450 ( .A(n163), .B(n155), .C(n156), .Q(n154) );
  OAI212 U468 ( .A(n185), .B(n195), .C(n186), .Q(n184) );
  XOR22 U507 ( .A(n33), .B(n262), .Q(SUM[5]) );
  AOI212 U515 ( .A(n588), .B(n548), .C(n473), .Q(n257) );
  XNR22 U516 ( .A(n25), .B(n207), .Q(SUM[13]) );
  OAI212 U517 ( .A(n208), .B(n584), .C(n209), .Q(n207) );
  XNR22 U518 ( .A(n12), .B(n90), .Q(SUM[26]) );
  OAI212 U527 ( .A(n599), .B(n566), .C(n602), .Q(n108) );
  OAI212 U529 ( .A(n188), .B(n584), .C(n189), .Q(n187) );
  OAI212 U533 ( .A(n244), .B(n584), .C(n564), .Q(n243) );
  OAI212 U539 ( .A(n256), .B(n252), .C(n253), .Q(n251) );
  XNR22 U540 ( .A(n10), .B(n72), .Q(SUM[28]) );
  XNR22 U542 ( .A(n24), .B(n196), .Q(SUM[14]) );
  XNR22 U550 ( .A(n9), .B(n63), .Q(SUM[29]) );
  XNR22 U557 ( .A(n11), .B(n81), .Q(SUM[27]) );
  XNR22 U561 ( .A(n31), .B(n254), .Q(SUM[7]) );
  XNR22 U562 ( .A(n14), .B(n108), .Q(SUM[24]) );
  XNR22 U574 ( .A(n23), .B(n187), .Q(SUM[15]) );
  OAI212 U663 ( .A(n241), .B(n564), .C(n242), .Q(n240) );
  NAND28 U398 ( .A(n448), .B(n449), .Q(SUM[21]) );
  OAI212 U349 ( .A(n53), .B(n550), .C(n54), .Q(n52) );
  BUF6 U350 ( .A(n258), .Q(n548) );
  CLKIN3 U351 ( .A(n566), .Q(n549) );
  INV6 U352 ( .A(n549), .Q(n550) );
  CLKIN4 U353 ( .A(n175), .Q(n570) );
  NAND22 U355 ( .A(n568), .B(n190), .Q(n188) );
  NAND24 U356 ( .A(n135), .B(n115), .Q(n113) );
  INV6 U357 ( .A(n247), .Q(n584) );
  OAI211 U358 ( .A(n597), .B(n566), .C(n600), .Q(n551) );
  NOR23 U359 ( .A(A[13]), .B(B[13]), .Q(n205) );
  OAI211 U360 ( .A(n194), .B(n625), .C(n195), .Q(n191) );
  INV2 U361 ( .A(n472), .Q(n625) );
  CLKIN6 U362 ( .A(n450), .Q(n575) );
  NAND24 U363 ( .A(n575), .B(n607), .Q(n471) );
  NAND22 U364 ( .A(A[3]), .B(B[3]), .Q(n272) );
  NOR23 U365 ( .A(B[3]), .B(A[3]), .Q(n271) );
  NOR24 U366 ( .A(A[6]), .B(B[6]), .Q(n255) );
  NAND23 U367 ( .A(A[6]), .B(B[6]), .Q(n256) );
  NAND28 U368 ( .A(n424), .B(n425), .Q(SUM[19]) );
  CLKIN3 U369 ( .A(n106), .Q(n641) );
  NOR23 U370 ( .A(n99), .B(n106), .Q(n97) );
  NAND24 U371 ( .A(n258), .B(n250), .Q(n248) );
  INV0 U372 ( .A(n260), .Q(n586) );
  NAND22 U373 ( .A(n157), .B(n19), .Q(n424) );
  CLKIN4 U374 ( .A(n157), .Q(n569) );
  NOR24 U375 ( .A(A[9]), .B(B[9]), .Q(n241) );
  NAND24 U376 ( .A(n436), .B(n437), .Q(SUM[25]) );
  OAI211 U377 ( .A(n213), .B(n205), .C(n206), .Q(n472) );
  NAND22 U378 ( .A(A[13]), .B(B[13]), .Q(n206) );
  NOR24 U380 ( .A(n117), .B(n126), .Q(n115) );
  NOR22 U381 ( .A(B[27]), .B(A[27]), .Q(n79) );
  XNR22 U382 ( .A(n26), .B(n214), .Q(SUM[12]) );
  XNR22 U383 ( .A(n28), .B(n232), .Q(SUM[10]) );
  NOR23 U384 ( .A(n255), .B(n252), .Q(n250) );
  INV3 U385 ( .A(n463), .Q(n601) );
  NAND24 U386 ( .A(n239), .B(n221), .Q(n219) );
  CLKIN6 U387 ( .A(n553), .Q(n554) );
  AOI210 U388 ( .A(n438), .B(n567), .C(n577), .Q(n227) );
  NOR22 U389 ( .A(B[16]), .B(A[16]), .Q(n176) );
  NAND22 U390 ( .A(n97), .B(n77), .Q(n6) );
  NOR21 U392 ( .A(n636), .B(n6), .Q(n55) );
  NOR23 U393 ( .A(A[11]), .B(B[11]), .Q(n223) );
  NOR22 U394 ( .A(A[21]), .B(B[21]), .Q(n137) );
  NOR21 U395 ( .A(n194), .B(n627), .Q(n190) );
  INV3 U396 ( .A(n135), .Q(n621) );
  AOI211 U397 ( .A(n204), .B(n183), .C(n184), .Q(n182) );
  NAND23 U399 ( .A(n203), .B(n183), .Q(n181) );
  NOR22 U400 ( .A(n113), .B(n151), .Q(n565) );
  NOR22 U401 ( .A(n70), .B(n6), .Q(n66) );
  AOI211 U402 ( .A(n576), .B(n632), .C(n631), .Q(n209) );
  AOI211 U403 ( .A(n601), .B(n624), .C(n622), .Q(n141) );
  CLKIN3 U404 ( .A(n139), .Q(n572) );
  CLKIN3 U405 ( .A(n243), .Q(n579) );
  INV3 U406 ( .A(n98), .Q(n612) );
  INV3 U407 ( .A(n119), .Q(n560) );
  NAND26 U408 ( .A(n461), .B(n462), .Q(SUM[20]) );
  NOR23 U409 ( .A(B[5]), .B(A[5]), .Q(n260) );
  NAND22 U410 ( .A(n470), .B(n471), .Q(SUM[18]) );
  NAND22 U411 ( .A(n551), .B(n20), .Q(n470) );
  INV3 U412 ( .A(n20), .Q(n607) );
  NAND24 U413 ( .A(n557), .B(n558), .Q(SUM[11]) );
  NAND23 U414 ( .A(n555), .B(n556), .Q(n558) );
  NAND22 U415 ( .A(n611), .B(n571), .Q(n437) );
  NAND26 U416 ( .A(n418), .B(n419), .Q(SUM[17]) );
  NAND24 U417 ( .A(n570), .B(n595), .Q(n419) );
  XOR21 U418 ( .A(n30), .B(n584), .Q(SUM[8]) );
  XOR21 U419 ( .A(n32), .B(n257), .Q(SUM[6]) );
  XNR21 U420 ( .A(n35), .B(n273), .Q(SUM[3]) );
  XOR21 U421 ( .A(n281), .B(n37), .Q(SUM[1]) );
  NAND26 U422 ( .A(n569), .B(n629), .Q(n425) );
  NOR24 U423 ( .A(B[7]), .B(A[7]), .Q(n252) );
  NAND22 U424 ( .A(B[5]), .B(A[5]), .Q(n261) );
  INV3 U425 ( .A(n112), .Q(n553) );
  OAI212 U426 ( .A(n597), .B(n566), .C(n600), .Q(n450) );
  CLKBU12 U427 ( .A(n566), .Q(n552) );
  OAI210 U428 ( .A(n266), .B(n260), .C(n261), .Q(n473) );
  CLKIN4 U429 ( .A(n146), .Q(n573) );
  NAND24 U430 ( .A(n171), .B(n153), .Q(n151) );
  NOR22 U431 ( .A(n173), .B(n176), .Q(n171) );
  NAND24 U432 ( .A(n561), .B(n562), .Q(SUM[23]) );
  NOR23 U434 ( .A(n155), .B(n162), .Q(n153) );
  NAND21 U435 ( .A(B[11]), .B(A[11]), .Q(n224) );
  NAND20 U436 ( .A(n617), .B(n118), .Q(n15) );
  NAND24 U437 ( .A(n623), .B(n573), .Q(n462) );
  NAND21 U438 ( .A(A[24]), .B(B[24]), .Q(n107) );
  NOR20 U439 ( .A(n444), .B(n274), .Q(n269) );
  XOR21 U440 ( .A(n36), .B(n594), .Q(SUM[2]) );
  OAI210 U441 ( .A(n274), .B(n594), .C(n275), .Q(n273) );
  NAND22 U442 ( .A(n225), .B(n27), .Q(n557) );
  INV3 U443 ( .A(n225), .Q(n555) );
  INV3 U444 ( .A(n27), .Q(n556) );
  BUF12 U445 ( .A(n245), .Q(n564) );
  INV0 U446 ( .A(n252), .Q(n585) );
  INV3 U447 ( .A(n101), .Q(n571) );
  INV1 U448 ( .A(n5), .Q(n613) );
  NOR22 U449 ( .A(B[22]), .B(A[22]), .Q(n126) );
  OAI210 U451 ( .A(n564), .B(n241), .C(n242), .Q(n438) );
  INV1 U452 ( .A(n438), .Q(n578) );
  CLKIN0 U453 ( .A(n241), .Q(n583) );
  NOR24 U454 ( .A(n185), .B(n194), .Q(n183) );
  NOR23 U455 ( .A(A[15]), .B(B[15]), .Q(n185) );
  NAND21 U456 ( .A(n608), .B(n163), .Q(n20) );
  NOR23 U457 ( .A(n181), .B(n219), .Q(n179) );
  NOR20 U458 ( .A(B[0]), .B(A[0]), .Q(n280) );
  AOI210 U459 ( .A(n554), .B(n66), .C(n67), .Q(n65) );
  NAND21 U460 ( .A(B[22]), .B(A[22]), .Q(n127) );
  NOR23 U461 ( .A(B[14]), .B(A[14]), .Q(n194) );
  NAND22 U462 ( .A(n15), .B(n119), .Q(n561) );
  NAND24 U463 ( .A(n559), .B(n560), .Q(n562) );
  INV3 U464 ( .A(n15), .Q(n559) );
  OAI212 U465 ( .A(n64), .B(n550), .C(n65), .Q(n63) );
  AOI211 U466 ( .A(n576), .B(n203), .C(n472), .Q(n198) );
  NOR23 U467 ( .A(B[12]), .B(A[12]), .Q(n212) );
  INV1 U469 ( .A(n576), .Q(n563) );
  NAND22 U470 ( .A(n605), .B(n256), .Q(n32) );
  NAND24 U471 ( .A(n582), .B(n579), .Q(n431) );
  NAND28 U472 ( .A(n430), .B(n431), .Q(SUM[9]) );
  AOI210 U473 ( .A(n554), .B(n616), .C(n613), .Q(n74) );
  NAND20 U474 ( .A(A[23]), .B(B[23]), .Q(n118) );
  NAND20 U475 ( .A(A[1]), .B(B[1]), .Q(n279) );
  NAND23 U476 ( .A(n139), .B(n17), .Q(n448) );
  NAND22 U477 ( .A(n29), .B(n243), .Q(n430) );
  NOR22 U478 ( .A(B[10]), .B(A[10]), .Q(n230) );
  OAI212 U479 ( .A(n73), .B(n552), .C(n74), .Q(n72) );
  AOI211 U480 ( .A(n554), .B(n84), .C(n85), .Q(n83) );
  NOR23 U481 ( .A(n223), .B(n230), .Q(n221) );
  NAND22 U482 ( .A(A[8]), .B(B[8]), .Q(n245) );
  NOR22 U483 ( .A(B[26]), .B(A[26]), .Q(n88) );
  NAND22 U484 ( .A(A[26]), .B(B[26]), .Q(n89) );
  INV2 U485 ( .A(n230), .Q(n567) );
  NOR23 U486 ( .A(n137), .B(n144), .Q(n135) );
  INV0 U487 ( .A(n126), .Q(n644) );
  INV0 U488 ( .A(n99), .Q(n614) );
  NOR22 U490 ( .A(B[25]), .B(A[25]), .Q(n99) );
  NOR21 U491 ( .A(n61), .B(n70), .Q(n59) );
  OAI211 U492 ( .A(n71), .B(n61), .C(n62), .Q(n60) );
  NOR21 U493 ( .A(B[29]), .B(A[29]), .Q(n61) );
  NAND20 U494 ( .A(n565), .B(n44), .Q(n42) );
  AOI211 U495 ( .A(n172), .B(n153), .C(n154), .Q(n463) );
  NAND22 U496 ( .A(A[20]), .B(B[20]), .Q(n145) );
  NAND21 U497 ( .A(A[21]), .B(B[21]), .Q(n138) );
  NOR22 U498 ( .A(B[20]), .B(A[20]), .Q(n144) );
  BUF15 U499 ( .A(n178), .Q(n566) );
  OAI211 U501 ( .A(n89), .B(n79), .C(n80), .Q(n78) );
  OAI212 U502 ( .A(n88), .B(n612), .C(n89), .Q(n85) );
  INV2 U503 ( .A(n220), .Q(n576) );
  OAI212 U504 ( .A(n220), .B(n181), .C(n182), .Q(n180) );
  AOI211 U505 ( .A(n601), .B(n135), .C(n136), .Q(n130) );
  NAND21 U506 ( .A(n598), .B(n135), .Q(n129) );
  NOR23 U508 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NAND20 U509 ( .A(n624), .B(n145), .Q(n18) );
  NAND22 U510 ( .A(n598), .B(n624), .Q(n140) );
  INV1 U511 ( .A(n144), .Q(n624) );
  AOI211 U513 ( .A(n554), .B(n97), .C(n98), .Q(n92) );
  NOR22 U514 ( .A(B[23]), .B(A[23]), .Q(n117) );
  NOR21 U519 ( .A(B[24]), .B(A[24]), .Q(n106) );
  NOR21 U520 ( .A(n88), .B(n615), .Q(n84) );
  INV0 U521 ( .A(n88), .Q(n640) );
  OAI211 U522 ( .A(n636), .B(n5), .C(n637), .Q(n56) );
  OAI211 U523 ( .A(n46), .B(n5), .C(n47), .Q(n45) );
  NOR22 U524 ( .A(n260), .B(n265), .Q(n258) );
  NOR22 U525 ( .A(B[17]), .B(A[17]), .Q(n173) );
  INV2 U526 ( .A(n212), .Q(n632) );
  CLKIN3 U528 ( .A(n79), .Q(n639) );
  NOR22 U530 ( .A(B[4]), .B(A[4]), .Q(n265) );
  INV1 U531 ( .A(n176), .Q(n609) );
  NOR22 U532 ( .A(n79), .B(n88), .Q(n77) );
  OAI211 U534 ( .A(n70), .B(n5), .C(n71), .Q(n67) );
  AOI212 U535 ( .A(n98), .B(n77), .C(n78), .Q(n5) );
  NAND22 U536 ( .A(n565), .B(n55), .Q(n53) );
  INV3 U537 ( .A(n219), .Q(n568) );
  NAND21 U538 ( .A(n568), .B(n203), .Q(n197) );
  NAND22 U541 ( .A(n565), .B(n66), .Q(n64) );
  NAND20 U543 ( .A(n583), .B(n242), .Q(n29) );
  NOR21 U544 ( .A(n113), .B(n151), .Q(n111) );
  NAND21 U545 ( .A(n272), .B(n587), .Q(n35) );
  INV3 U546 ( .A(n151), .Q(n598) );
  CLKIN0 U547 ( .A(n136), .Q(n619) );
  NOR21 U548 ( .A(n126), .B(n621), .Q(n122) );
  OAI211 U549 ( .A(n126), .B(n619), .C(n127), .Q(n123) );
  NAND21 U551 ( .A(n16), .B(n128), .Q(n455) );
  NAND26 U552 ( .A(n572), .B(n618), .Q(n449) );
  CLKIN3 U553 ( .A(n97), .Q(n615) );
  NAND20 U554 ( .A(n641), .B(n107), .Q(n14) );
  CLKIN3 U555 ( .A(n111), .Q(n599) );
  INV0 U556 ( .A(n162), .Q(n608) );
  NAND21 U558 ( .A(n565), .B(n616), .Q(n73) );
  NAND21 U559 ( .A(n111), .B(n97), .Q(n91) );
  XNR21 U560 ( .A(n34), .B(n588), .Q(SUM[4]) );
  INV0 U563 ( .A(n255), .Q(n605) );
  NOR20 U564 ( .A(n46), .B(n6), .Q(n44) );
  NAND21 U565 ( .A(n568), .B(n632), .Q(n208) );
  INV0 U566 ( .A(n231), .Q(n577) );
  NAND24 U567 ( .A(n455), .B(n456), .Q(SUM[22]) );
  NAND22 U568 ( .A(n643), .B(n574), .Q(n456) );
  NAND20 U569 ( .A(n596), .B(n174), .Q(n21) );
  NAND20 U570 ( .A(n644), .B(n127), .Q(n16) );
  INV0 U571 ( .A(n194), .Q(n610) );
  NAND20 U572 ( .A(n171), .B(n608), .Q(n158) );
  NAND20 U573 ( .A(A[28]), .B(B[28]), .Q(n71) );
  NAND20 U575 ( .A(A[31]), .B(B[31]), .Q(n40) );
  NAND20 U576 ( .A(A[30]), .B(B[30]), .Q(n51) );
  NAND20 U577 ( .A(A[27]), .B(B[27]), .Q(n80) );
  INV3 U578 ( .A(n29), .Q(n582) );
  INV3 U579 ( .A(n128), .Q(n574) );
  NAND20 U580 ( .A(n239), .B(n567), .Q(n226) );
  INV3 U581 ( .A(n6), .Q(n616) );
  NAND20 U582 ( .A(n261), .B(n586), .Q(n33) );
  NAND20 U583 ( .A(n609), .B(n177), .Q(n22) );
  NAND22 U584 ( .A(n580), .B(n564), .Q(n30) );
  INV0 U585 ( .A(n244), .Q(n580) );
  NAND20 U586 ( .A(n589), .B(n266), .Q(n34) );
  NAND20 U587 ( .A(n585), .B(n253), .Q(n31) );
  CLKIN0 U588 ( .A(n239), .Q(n581) );
  INV3 U589 ( .A(n60), .Q(n637) );
  INV0 U590 ( .A(n205), .Q(n626) );
  NAND20 U591 ( .A(n604), .B(n224), .Q(n27) );
  NAND22 U592 ( .A(n175), .B(n21), .Q(n418) );
  INV3 U593 ( .A(n21), .Q(n595) );
  INV3 U594 ( .A(n19), .Q(n629) );
  NAND21 U595 ( .A(n111), .B(n84), .Q(n82) );
  NAND22 U596 ( .A(n18), .B(n146), .Q(n461) );
  INV3 U597 ( .A(n18), .Q(n623) );
  INV3 U598 ( .A(n16), .Q(n643) );
  NAND22 U599 ( .A(n101), .B(n13), .Q(n436) );
  INV3 U600 ( .A(n13), .Q(n611) );
  INV3 U601 ( .A(n17), .Q(n618) );
  CLKIN0 U602 ( .A(n172), .Q(n600) );
  NAND22 U603 ( .A(n598), .B(n122), .Q(n120) );
  INV0 U604 ( .A(n266), .Q(n590) );
  INV3 U605 ( .A(n59), .Q(n636) );
  INV3 U606 ( .A(n265), .Q(n589) );
  INV3 U607 ( .A(n171), .Q(n597) );
  INV3 U608 ( .A(n277), .Q(n594) );
  NAND20 U609 ( .A(n591), .B(n275), .Q(n36) );
  INV2 U610 ( .A(n274), .Q(n591) );
  NAND20 U611 ( .A(n186), .B(n603), .Q(n23) );
  INV0 U612 ( .A(n185), .Q(n603) );
  NAND20 U613 ( .A(n610), .B(n195), .Q(n24) );
  INV2 U614 ( .A(n444), .Q(n587) );
  AOI210 U615 ( .A(n172), .B(n608), .C(n606), .Q(n159) );
  INV0 U616 ( .A(n163), .Q(n606) );
  NAND22 U617 ( .A(n634), .B(n51), .Q(n8) );
  INV0 U618 ( .A(n117), .Q(n617) );
  NAND22 U619 ( .A(n638), .B(n62), .Q(n9) );
  INV3 U620 ( .A(n61), .Q(n638) );
  AOI210 U621 ( .A(n60), .B(n634), .C(n633), .Q(n47) );
  INV3 U622 ( .A(n51), .Q(n633) );
  INV3 U623 ( .A(n145), .Q(n622) );
  NAND22 U624 ( .A(n635), .B(n71), .Q(n10) );
  INV0 U625 ( .A(n70), .Q(n635) );
  NAND22 U626 ( .A(n640), .B(n89), .Q(n12) );
  NAND22 U627 ( .A(n639), .B(n80), .Q(n11) );
  NAND22 U628 ( .A(n628), .B(n279), .Q(n37) );
  INV2 U629 ( .A(n278), .Q(n628) );
  NAND22 U630 ( .A(n565), .B(n641), .Q(n102) );
  INV3 U631 ( .A(n107), .Q(n642) );
  NAND21 U632 ( .A(n630), .B(n156), .Q(n19) );
  INV0 U633 ( .A(n155), .Q(n630) );
  INV0 U634 ( .A(n173), .Q(n596) );
  NAND20 U635 ( .A(n614), .B(n100), .Q(n13) );
  AOI211 U636 ( .A(n601), .B(n122), .C(n123), .Q(n121) );
  INV0 U637 ( .A(n213), .Q(n631) );
  NAND21 U638 ( .A(n620), .B(n138), .Q(n17) );
  INV0 U639 ( .A(n137), .Q(n620) );
  NAND21 U640 ( .A(n59), .B(n634), .Q(n46) );
  XNR21 U641 ( .A(n7), .B(n41), .Q(SUM[31]) );
  NAND22 U642 ( .A(n645), .B(n40), .Q(n7) );
  NAND20 U643 ( .A(A[29]), .B(B[29]), .Q(n62) );
  INV3 U644 ( .A(n50), .Q(n634) );
  NOR20 U645 ( .A(B[30]), .B(A[30]), .Q(n50) );
  INV3 U646 ( .A(n38), .Q(SUM[0]) );
  NAND22 U647 ( .A(n593), .B(n281), .Q(n38) );
  INV3 U648 ( .A(n280), .Q(n593) );
  INV3 U649 ( .A(n39), .Q(n645) );
  NOR20 U650 ( .A(B[31]), .B(A[31]), .Q(n39) );
  NAND20 U651 ( .A(A[0]), .B(B[0]), .Q(n281) );
  NAND21 U652 ( .A(A[19]), .B(B[19]), .Q(n156) );
  NAND21 U653 ( .A(A[25]), .B(B[25]), .Q(n100) );
  NOR21 U654 ( .A(B[2]), .B(A[2]), .Q(n274) );
  NAND21 U655 ( .A(n567), .B(n231), .Q(n28) );
  NAND22 U656 ( .A(A[10]), .B(B[10]), .Q(n231) );
  OAI211 U657 ( .A(n213), .B(n205), .C(n206), .Q(n204) );
  NAND21 U658 ( .A(n626), .B(n206), .Q(n25) );
  OAI212 U659 ( .A(n275), .B(n271), .C(n272), .Q(n270) );
  NAND22 U660 ( .A(n632), .B(n213), .Q(n26) );
  INV2 U661 ( .A(n223), .Q(n604) );
  OAI212 U662 ( .A(n255), .B(n257), .C(n256), .Q(n254) );
  OAI212 U664 ( .A(n266), .B(n260), .C(n261), .Q(n259) );
  INV1 U665 ( .A(n203), .Q(n627) );
  NOR22 U666 ( .A(B[28]), .B(A[28]), .Q(n70) );
  AOI211 U667 ( .A(n576), .B(n190), .C(n191), .Q(n189) );
  XNR22 U668 ( .A(n8), .B(n52), .Q(SUM[30]) );
  NOR23 U669 ( .A(n241), .B(n244), .Q(n239) );
  NOR20 U670 ( .A(B[1]), .B(A[1]), .Q(n278) );
  OAI212 U671 ( .A(n82), .B(n566), .C(n83), .Q(n81) );
  NAND21 U672 ( .A(B[15]), .B(A[15]), .Q(n186) );
  NAND21 U673 ( .A(A[17]), .B(B[17]), .Q(n174) );
  NOR22 U674 ( .A(B[18]), .B(A[18]), .Q(n162) );
  NAND22 U675 ( .A(A[18]), .B(B[18]), .Q(n163) );
  OAI212 U676 ( .A(n102), .B(n566), .C(n103), .Q(n101) );
  AOI211 U677 ( .A(n112), .B(n641), .C(n642), .Q(n103) );
  NAND22 U678 ( .A(B[14]), .B(A[14]), .Q(n195) );
  NAND22 U679 ( .A(A[12]), .B(B[12]), .Q(n213) );
  NAND21 U680 ( .A(A[7]), .B(B[7]), .Q(n253) );
  NAND22 U681 ( .A(A[16]), .B(B[16]), .Q(n177) );
  NAND23 U682 ( .A(A[4]), .B(B[4]), .Q(n266) );
  NAND23 U683 ( .A(B[2]), .B(A[2]), .Q(n275) );
  OAI210 U684 ( .A(n42), .B(n552), .C(n43), .Q(n41) );
  INV2 U685 ( .A(n268), .Q(n588) );
  NAND22 U686 ( .A(B[9]), .B(A[9]), .Q(n242) );
  OAI211 U687 ( .A(n219), .B(n584), .C(n563), .Q(n214) );
  INV1 U688 ( .A(n554), .Q(n602) );
  NOR20 U689 ( .A(A[3]), .B(B[3]), .Q(n444) );
  NOR22 U690 ( .A(B[8]), .B(A[8]), .Q(n244) );
  AOI210 U691 ( .A(n554), .B(n44), .C(n45), .Q(n43) );
  AOI210 U692 ( .A(n554), .B(n55), .C(n56), .Q(n54) );
endmodule


module adder_1 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   n1;

  adder_1_DW01_add_1 add_16 ( .A(A), .B(B), .CI(n1), .SUM(O) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module iir_sol ( Reset, Clk, Input, Output );
  input [319:0] Input;
  output [31:0] Output;
  input Reset, Clk;
  wire   s_80__31_, s_80__30_, s_80__29_, s_80__28_, s_80__27_, s_80__26_,
         s_80__25_, s_80__24_, s_80__23_, s_80__22_, s_80__21_, s_80__20_,
         s_80__19_, s_80__18_, s_80__17_, s_80__16_, s_80__15_, s_80__14_,
         s_80__13_, s_80__12_, s_80__11_, s_80__10_, s_80__9_, s_80__8_,
         s_80__7_, s_80__6_, s_80__5_, s_80__4_, s_80__3_, s_80__2_, s_80__1_,
         s_80__0_, s_81__31_, s_81__30_, s_81__29_, s_81__28_, s_81__27_,
         s_81__26_, s_81__25_, s_81__24_, s_81__23_, s_81__22_, s_81__21_,
         s_81__20_, s_81__19_, s_81__18_, s_81__17_, s_81__16_, s_81__15_,
         s_81__14_, s_81__13_, s_81__12_, s_81__11_, s_81__10_, s_81__9_,
         s_81__8_, s_81__7_, s_81__6_, s_81__5_, s_81__4_, s_81__3_, s_81__2_,
         s_81__1_, s_81__0_, s_82__31_, s_82__30_, s_82__29_, s_82__28_,
         s_82__27_, s_82__26_, s_82__25_, s_82__24_, s_82__23_, s_82__22_,
         s_82__21_, s_82__20_, s_82__19_, s_82__18_, s_82__17_, s_82__16_,
         s_82__15_, s_82__14_, s_82__13_, s_82__12_, s_82__11_, s_82__10_,
         s_82__9_, s_82__8_, s_82__7_, s_82__6_, s_82__5_, s_82__4_, s_82__3_,
         s_82__2_, s_82__1_, s_82__0_, s_83__31_, s_83__30_, s_83__29_,
         s_83__28_, s_83__27_, s_83__26_, s_83__25_, s_83__24_, s_83__23_,
         s_83__22_, s_83__21_, s_83__20_, s_83__19_, s_83__18_, s_83__17_,
         s_83__16_, s_83__15_, s_83__14_, s_83__13_, s_83__12_, s_83__11_,
         s_83__10_, s_83__9_, s_83__8_, s_83__7_, s_83__6_, s_83__5_, s_83__4_,
         s_83__3_, s_83__2_, s_83__1_, s_83__0_, s_84__31_, s_84__30_,
         s_84__29_, s_84__28_, s_84__27_, s_84__26_, s_84__25_, s_84__24_,
         s_84__23_, s_84__22_, s_84__21_, s_84__20_, s_84__19_, s_84__18_,
         s_84__17_, s_84__16_, s_84__15_, s_84__14_, s_84__13_, s_84__12_,
         s_84__11_, s_84__10_, s_84__9_, s_84__8_, s_84__7_, s_84__6_,
         s_84__5_, s_84__4_, s_84__3_, s_84__2_, s_84__1_, s_84__0_, s_85__31_,
         s_85__30_, s_85__29_, s_85__28_, s_85__27_, s_85__26_, s_85__25_,
         s_85__24_, s_85__23_, s_85__22_, s_85__21_, s_85__20_, s_85__19_,
         s_85__18_, s_85__17_, s_85__16_, s_85__15_, s_85__14_, s_85__13_,
         s_85__12_, s_85__11_, s_85__10_, s_85__9_, s_85__8_, s_85__7_,
         s_85__6_, s_85__5_, s_85__4_, s_85__3_, s_85__2_, s_85__1_, s_85__0_,
         s_86__31_, s_86__30_, s_86__29_, s_86__28_, s_86__27_, s_86__26_,
         s_86__25_, s_86__24_, s_86__23_, s_86__22_, s_86__21_, s_86__20_,
         s_86__19_, s_86__18_, s_86__17_, s_86__16_, s_86__15_, s_86__14_,
         s_86__13_, s_86__12_, s_86__11_, s_86__10_, s_86__9_, s_86__8_,
         s_86__7_, s_86__6_, s_86__5_, s_86__4_, s_86__3_, s_86__2_, s_86__1_,
         s_86__0_, s_87__31_, s_87__30_, s_87__29_, s_87__28_, s_87__27_,
         s_87__26_, s_87__25_, s_87__24_, s_87__23_, s_87__22_, s_87__21_,
         s_87__20_, s_87__19_, s_87__18_, s_87__17_, s_87__16_, s_87__15_,
         s_87__14_, s_87__13_, s_87__12_, s_87__11_, s_87__10_, s_87__9_,
         s_87__8_, s_87__7_, s_87__6_, s_87__5_, s_87__4_, s_87__3_, s_87__2_,
         s_87__1_, s_87__0_, s_88__31_, s_88__30_, s_88__29_, s_88__28_,
         s_88__27_, s_88__26_, s_88__25_, s_88__24_, s_88__23_, s_88__22_,
         s_88__21_, s_88__20_, s_88__19_, s_88__18_, s_88__17_, s_88__16_,
         s_88__15_, s_88__14_, s_88__13_, s_88__12_, s_88__11_, s_88__10_,
         s_88__9_, s_88__8_, s_88__7_, s_88__6_, s_88__5_, s_88__4_, s_88__3_,
         s_88__2_, s_88__1_, s_88__0_, s_89__31_, s_89__30_, s_89__29_,
         s_89__28_, s_89__27_, s_89__26_, s_89__25_, s_89__24_, s_89__23_,
         s_89__22_, s_89__21_, s_89__20_, s_89__19_, s_89__18_, s_89__17_,
         s_89__16_, s_89__15_, s_89__14_, s_89__13_, s_89__12_, s_89__11_,
         s_89__10_, s_89__9_, s_89__8_, s_89__7_, s_89__6_, s_89__5_, s_89__4_,
         s_89__3_, s_89__2_, s_89__1_, s_89__0_, s_90__31_, s_90__30_,
         s_90__29_, s_90__28_, s_90__27_, s_90__26_, s_90__25_, s_90__24_,
         s_90__23_, s_90__22_, s_90__21_, s_90__20_, s_90__19_, s_90__18_,
         s_90__17_, s_90__16_, s_90__15_, s_90__14_, s_90__13_, s_90__12_,
         s_90__11_, s_90__10_, s_90__9_, s_90__8_, s_90__7_, s_90__6_,
         s_90__5_, s_90__4_, s_90__3_, s_90__2_, s_90__1_, s_90__0_, s_91__31_,
         s_91__30_, s_91__29_, s_91__28_, s_91__27_, s_91__26_, s_91__25_,
         s_91__24_, s_91__23_, s_91__22_, s_91__21_, s_91__20_, s_91__19_,
         s_91__18_, s_91__17_, s_91__16_, s_91__15_, s_91__14_, s_91__13_,
         s_91__12_, s_91__11_, s_91__10_, s_91__9_, s_91__8_, s_91__7_,
         s_91__6_, s_91__5_, s_91__4_, s_91__3_, s_91__2_, s_91__1_, s_91__0_,
         y_1__31_, y_1__30_, y_1__29_, y_1__28_, y_1__27_, y_1__26_, y_1__25_,
         y_1__24_, y_1__23_, y_1__22_, y_1__21_, y_1__20_, y_1__19_, y_1__18_,
         y_1__17_, y_1__16_, y_1__15_, y_1__14_, y_1__13_, y_1__12_, y_1__11_,
         y_1__10_, y_1__9_, y_1__8_, y_1__7_, y_1__6_, y_1__5_, y_1__4_,
         y_1__3_, y_1__2_, y_1__1_, y_1__0_, y_2__31_, y_2__30_, y_2__29_,
         y_2__28_, y_2__27_, y_2__26_, y_2__25_, y_2__24_, y_2__23_, y_2__22_,
         y_2__21_, y_2__20_, y_2__19_, y_2__18_, y_2__17_, y_2__16_, y_2__15_,
         y_2__14_, y_2__13_, y_2__12_, y_2__11_, y_2__10_, y_2__9_, y_2__8_,
         y_2__7_, y_2__6_, y_2__5_, y_2__4_, y_2__3_, y_2__2_, y_2__1_,
         y_2__0_, y_3__31_, y_3__30_, y_3__29_, y_3__28_, y_3__27_, y_3__26_,
         y_3__25_, y_3__24_, y_3__23_, y_3__22_, y_3__21_, y_3__20_, y_3__19_,
         y_3__18_, y_3__17_, y_3__16_, y_3__15_, y_3__14_, y_3__13_, y_3__12_,
         y_3__11_, y_3__10_, y_3__9_, y_3__8_, y_3__7_, y_3__6_, y_3__5_,
         y_3__4_, y_3__3_, y_3__2_, y_3__1_, y_3__0_, y_4__31_, y_4__30_,
         y_4__29_, y_4__28_, y_4__27_, y_4__26_, y_4__25_, y_4__24_, y_4__23_,
         y_4__22_, y_4__21_, y_4__20_, y_4__19_, y_4__18_, y_4__17_, y_4__16_,
         y_4__15_, y_4__14_, y_4__13_, y_4__12_, y_4__11_, y_4__10_, y_4__9_,
         y_4__8_, y_4__7_, y_4__6_, y_4__5_, y_4__4_, y_4__3_, y_4__2_,
         y_4__1_, y_4__0_, y_5__31_, y_5__30_, y_5__29_, y_5__28_, y_5__27_,
         y_5__26_, y_5__25_, y_5__24_, y_5__23_, y_5__22_, y_5__21_, y_5__20_,
         y_5__19_, y_5__18_, y_5__17_, y_5__16_, y_5__15_, y_5__14_, y_5__13_,
         y_5__12_, y_5__11_, y_5__10_, y_5__9_, y_5__8_, y_5__7_, y_5__6_,
         y_5__5_, y_5__4_, y_5__3_, y_5__2_, y_5__1_, y_5__0_, y_6__31_,
         y_6__30_, y_6__29_, y_6__28_, y_6__27_, y_6__26_, y_6__25_, y_6__24_,
         y_6__23_, y_6__22_, y_6__21_, y_6__20_, y_6__19_, y_6__18_, y_6__17_,
         y_6__16_, y_6__15_, y_6__14_, y_6__13_, y_6__12_, y_6__11_, y_6__10_,
         y_6__9_, y_6__8_, y_6__7_, y_6__6_, y_6__5_, y_6__4_, y_6__3_,
         y_6__2_, y_6__1_, y_6__0_, y_7__31_, y_7__30_, y_7__29_, y_7__28_,
         y_7__27_, y_7__26_, y_7__25_, y_7__24_, y_7__23_, y_7__22_, y_7__21_,
         y_7__20_, y_7__19_, y_7__18_, y_7__17_, y_7__16_, y_7__15_, y_7__14_,
         y_7__13_, y_7__12_, y_7__11_, y_7__10_, y_7__9_, y_7__8_, y_7__7_,
         y_7__6_, y_7__5_, y_7__4_, y_7__3_, y_7__2_, y_7__1_, y_7__0_,
         y_8__31_, y_8__30_, y_8__29_, y_8__28_, y_8__27_, y_8__26_, y_8__25_,
         y_8__24_, y_8__23_, y_8__22_, y_8__21_, y_8__20_, y_8__19_, y_8__18_,
         y_8__17_, y_8__16_, y_8__15_, y_8__14_, y_8__13_, y_8__12_, y_8__11_,
         y_8__10_, y_8__9_, y_8__8_, y_8__7_, y_8__6_, y_8__5_, y_8__4_,
         y_8__3_, y_8__2_, y_8__1_, y_8__0_, s_47__31_, s_47__30_, s_47__29_,
         s_47__28_, s_47__27_, s_47__26_, s_47__25_, s_47__24_, s_47__23_,
         s_47__22_, s_47__21_, s_47__20_, s_47__19_, s_47__18_, s_47__17_,
         s_47__16_, s_47__15_, s_47__14_, s_47__13_, s_47__12_, s_47__11_,
         s_47__10_, s_47__9_, s_47__8_, s_47__7_, s_47__6_, s_47__5_, s_47__4_,
         s_47__3_, s_47__2_, s_47__1_, s_47__0_, s_48__31_, s_48__30_,
         s_48__29_, s_48__28_, s_48__27_, s_48__26_, s_48__25_, s_48__24_,
         s_48__23_, s_48__22_, s_48__21_, s_48__20_, s_48__19_, s_48__18_,
         s_48__17_, s_48__16_, s_48__15_, s_48__14_, s_48__13_, s_48__12_,
         s_48__11_, s_48__10_, s_48__9_, s_48__8_, s_48__7_, s_48__6_,
         s_48__5_, s_48__4_, s_48__3_, s_48__2_, s_48__1_, s_48__0_, s_49__31_,
         s_49__30_, s_49__29_, s_49__28_, s_49__27_, s_49__26_, s_49__25_,
         s_49__24_, s_49__23_, s_49__22_, s_49__21_, s_49__20_, s_49__19_,
         s_49__18_, s_49__17_, s_49__16_, s_49__15_, s_49__14_, s_49__13_,
         s_49__12_, s_49__11_, s_49__10_, s_49__9_, s_49__8_, s_49__7_,
         s_49__6_, s_49__5_, s_49__4_, s_49__3_, s_49__2_, s_49__1_, s_49__0_,
         s_50__31_, s_50__30_, s_50__29_, s_50__28_, s_50__27_, s_50__26_,
         s_50__25_, s_50__24_, s_50__23_, s_50__22_, s_50__21_, s_50__20_,
         s_50__19_, s_50__18_, s_50__17_, s_50__16_, s_50__15_, s_50__14_,
         s_50__13_, s_50__12_, s_50__11_, s_50__10_, s_50__9_, s_50__8_,
         s_50__7_, s_50__6_, s_50__5_, s_50__4_, s_50__3_, s_50__2_, s_50__1_,
         s_50__0_, s_51__31_, s_51__30_, s_51__29_, s_51__28_, s_51__27_,
         s_51__26_, s_51__25_, s_51__24_, s_51__23_, s_51__22_, s_51__21_,
         s_51__20_, s_51__19_, s_51__18_, s_51__17_, s_51__16_, s_51__15_,
         s_51__14_, s_51__13_, s_51__12_, s_51__11_, s_51__10_, s_51__9_,
         s_51__8_, s_51__7_, s_51__6_, s_51__5_, s_51__4_, s_51__3_, s_51__2_,
         s_51__1_, s_51__0_, s_52__31_, s_52__30_, s_52__29_, s_52__28_,
         s_52__27_, s_52__26_, s_52__25_, s_52__24_, s_52__23_, s_52__22_,
         s_52__21_, s_52__20_, s_52__19_, s_52__18_, s_52__17_, s_52__16_,
         s_52__15_, s_52__14_, s_52__13_, s_52__12_, s_52__11_, s_52__10_,
         s_52__9_, s_52__8_, s_52__7_, s_52__6_, s_52__5_, s_52__4_, s_52__3_,
         s_52__2_, s_52__1_, s_52__0_, s_53__31_, s_53__30_, s_53__29_,
         s_53__28_, s_53__27_, s_53__26_, s_53__25_, s_53__24_, s_53__23_,
         s_53__22_, s_53__21_, s_53__20_, s_53__19_, s_53__18_, s_53__17_,
         s_53__16_, s_53__15_, s_53__14_, s_53__13_, s_53__12_, s_53__11_,
         s_53__10_, s_53__9_, s_53__8_, s_53__7_, s_53__6_, s_53__5_, s_53__4_,
         s_53__3_, s_53__2_, s_53__1_, s_53__0_, s_54__31_, s_54__30_,
         s_54__29_, s_54__28_, s_54__27_, s_54__26_, s_54__25_, s_54__24_,
         s_54__23_, s_54__22_, s_54__21_, s_54__20_, s_54__19_, s_54__18_,
         s_54__17_, s_54__16_, s_54__15_, s_54__14_, s_54__13_, s_54__12_,
         s_54__11_, s_54__10_, s_54__9_, s_54__8_, s_54__7_, s_54__6_,
         s_54__5_, s_54__4_, s_54__3_, s_54__2_, s_54__1_, s_54__0_, s_55__31_,
         s_55__30_, s_55__29_, s_55__28_, s_55__27_, s_55__26_, s_55__25_,
         s_55__24_, s_55__23_, s_55__22_, s_55__21_, s_55__20_, s_55__19_,
         s_55__18_, s_55__17_, s_55__16_, s_55__15_, s_55__14_, s_55__13_,
         s_55__12_, s_55__11_, s_55__10_, s_55__9_, s_55__8_, s_55__7_,
         s_55__6_, s_55__5_, s_55__4_, s_55__3_, s_55__2_, s_55__1_, s_55__0_,
         s_56__31_, s_56__30_, s_56__29_, s_56__28_, s_56__27_, s_56__26_,
         s_56__25_, s_56__24_, s_56__23_, s_56__22_, s_56__21_, s_56__20_,
         s_56__19_, s_56__18_, s_56__17_, s_56__16_, s_56__15_, s_56__14_,
         s_56__13_, s_56__12_, s_56__11_, s_56__10_, s_56__9_, s_56__8_,
         s_56__7_, s_56__6_, s_56__5_, s_56__4_, s_56__3_, s_56__2_, s_56__1_,
         s_56__0_, s_57__31_, s_57__30_, s_57__29_, s_57__28_, s_57__27_,
         s_57__26_, s_57__25_, s_57__24_, s_57__23_, s_57__22_, s_57__21_,
         s_57__20_, s_57__19_, s_57__18_, s_57__17_, s_57__16_, s_57__15_,
         s_57__14_, s_57__13_, s_57__12_, s_57__11_, s_57__10_, s_57__9_,
         s_57__8_, s_57__7_, s_57__6_, s_57__5_, s_57__4_, s_57__3_, s_57__2_,
         s_57__1_, s_57__0_, s_58__31_, s_58__30_, s_58__29_, s_58__28_,
         s_58__27_, s_58__26_, s_58__25_, s_58__24_, s_58__23_, s_58__22_,
         s_58__21_, s_58__20_, s_58__19_, s_58__18_, s_58__17_, s_58__16_,
         s_58__15_, s_58__14_, s_58__13_, s_58__12_, s_58__11_, s_58__10_,
         s_58__9_, s_58__8_, s_58__7_, s_58__6_, s_58__5_, s_58__4_, s_58__3_,
         s_58__2_, s_58__1_, s_58__0_, s_59__31_, s_59__30_, s_59__29_,
         s_59__28_, s_59__27_, s_59__26_, s_59__25_, s_59__24_, s_59__23_,
         s_59__22_, s_59__21_, s_59__20_, s_59__19_, s_59__18_, s_59__17_,
         s_59__16_, s_59__15_, s_59__14_, s_59__13_, s_59__12_, s_59__11_,
         s_59__10_, s_59__9_, s_59__8_, s_59__7_, s_59__6_, s_59__5_, s_59__4_,
         s_59__3_, s_59__2_, s_59__1_, s_59__0_, s_60__31_, s_60__30_,
         s_60__29_, s_60__28_, s_60__27_, s_60__26_, s_60__25_, s_60__24_,
         s_60__23_, s_60__22_, s_60__21_, s_60__20_, s_60__19_, s_60__18_,
         s_60__17_, s_60__16_, s_60__15_, s_60__14_, s_60__13_, s_60__12_,
         s_60__11_, s_60__10_, s_60__9_, s_60__8_, s_60__7_, s_60__6_,
         s_60__5_, s_60__4_, s_60__3_, s_60__2_, s_60__1_, s_60__0_, s_61__31_,
         s_61__30_, s_61__29_, s_61__28_, s_61__27_, s_61__26_, s_61__25_,
         s_61__24_, s_61__23_, s_61__22_, s_61__21_, s_61__20_, s_61__19_,
         s_61__18_, s_61__17_, s_61__16_, s_61__15_, s_61__14_, s_61__13_,
         s_61__12_, s_61__11_, s_61__10_, s_61__9_, s_61__8_, s_61__7_,
         s_61__6_, s_61__5_, s_61__4_, s_61__3_, s_61__2_, s_61__1_, s_61__0_,
         s_62__31_, s_62__30_, s_62__29_, s_62__28_, s_62__27_, s_62__26_,
         s_62__25_, s_62__24_, s_62__23_, s_62__22_, s_62__21_, s_62__20_,
         s_62__19_, s_62__18_, s_62__17_, s_62__16_, s_62__15_, s_62__14_,
         s_62__13_, s_62__12_, s_62__11_, s_62__10_, s_62__9_, s_62__8_,
         s_62__7_, s_62__6_, s_62__5_, s_62__4_, s_62__3_, s_62__2_, s_62__1_,
         s_62__0_, s_63__31_, s_63__30_, s_63__29_, s_63__28_, s_63__27_,
         s_63__26_, s_63__25_, s_63__24_, s_63__23_, s_63__22_, s_63__21_,
         s_63__20_, s_63__19_, s_63__18_, s_63__17_, s_63__16_, s_63__15_,
         s_63__14_, s_63__13_, s_63__12_, s_63__11_, s_63__10_, s_63__9_,
         s_63__8_, s_63__7_, s_63__6_, s_63__5_, s_63__4_, s_63__3_, s_63__2_,
         s_63__1_, s_63__0_, s_64__31_, s_64__30_, s_64__29_, s_64__28_,
         s_64__27_, s_64__26_, s_64__25_, s_64__24_, s_64__23_, s_64__22_,
         s_64__21_, s_64__20_, s_64__19_, s_64__18_, s_64__17_, s_64__16_,
         s_64__15_, s_64__14_, s_64__13_, s_64__12_, s_64__11_, s_64__10_,
         s_64__9_, s_64__8_, s_64__7_, s_64__6_, s_64__5_, s_64__4_, s_64__3_,
         s_64__2_, s_64__1_, s_64__0_, s_65__31_, s_65__30_, s_65__29_,
         s_65__28_, s_65__27_, s_65__26_, s_65__25_, s_65__24_, s_65__23_,
         s_65__22_, s_65__21_, s_65__20_, s_65__19_, s_65__18_, s_65__17_,
         s_65__16_, s_65__15_, s_65__14_, s_65__13_, s_65__12_, s_65__11_,
         s_65__10_, s_65__9_, s_65__8_, s_65__7_, s_65__6_, s_65__5_, s_65__4_,
         s_65__3_, s_65__2_, s_65__1_, s_65__0_, s_66__31_, s_66__30_,
         s_66__29_, s_66__28_, s_66__27_, s_66__26_, s_66__25_, s_66__24_,
         s_66__23_, s_66__22_, s_66__21_, s_66__20_, s_66__19_, s_66__18_,
         s_66__17_, s_66__16_, s_66__15_, s_66__14_, s_66__13_, s_66__12_,
         s_66__11_, s_66__10_, s_66__9_, s_66__8_, s_66__7_, s_66__6_,
         s_66__5_, s_66__4_, s_66__3_, s_66__2_, s_66__1_, s_66__0_, s_67__31_,
         s_67__30_, s_67__29_, s_67__28_, s_67__27_, s_67__26_, s_67__25_,
         s_67__24_, s_67__23_, s_67__22_, s_67__21_, s_67__20_, s_67__19_,
         s_67__18_, s_67__17_, s_67__16_, s_67__15_, s_67__14_, s_67__13_,
         s_67__12_, s_67__11_, s_67__10_, s_67__9_, s_67__8_, s_67__7_,
         s_67__6_, s_67__5_, s_67__4_, s_67__3_, s_67__2_, s_67__1_, s_67__0_,
         s_68__31_, s_68__30_, s_68__29_, s_68__28_, s_68__27_, s_68__26_,
         s_68__25_, s_68__24_, s_68__23_, s_68__22_, s_68__21_, s_68__20_,
         s_68__19_, s_68__18_, s_68__17_, s_68__16_, s_68__15_, s_68__14_,
         s_68__13_, s_68__12_, s_68__11_, s_68__10_, s_68__9_, s_68__8_,
         s_68__7_, s_68__6_, s_68__5_, s_68__4_, s_68__3_, s_68__2_, s_68__1_,
         s_68__0_, s_69__31_, s_69__30_, s_69__29_, s_69__28_, s_69__27_,
         s_69__26_, s_69__25_, s_69__24_, s_69__23_, s_69__22_, s_69__21_,
         s_69__20_, s_69__19_, s_69__18_, s_69__17_, s_69__16_, s_69__15_,
         s_69__14_, s_69__13_, s_69__12_, s_69__11_, s_69__10_, s_69__9_,
         s_69__8_, s_69__7_, s_69__6_, s_69__5_, s_69__4_, s_69__3_, s_69__2_,
         s_69__1_, s_69__0_, s_70__31_, s_70__30_, s_70__29_, s_70__28_,
         s_70__27_, s_70__26_, s_70__25_, s_70__24_, s_70__23_, s_70__22_,
         s_70__21_, s_70__20_, s_70__19_, s_70__18_, s_70__17_, s_70__16_,
         s_70__15_, s_70__14_, s_70__13_, s_70__12_, s_70__11_, s_70__10_,
         s_70__9_, s_70__8_, s_70__7_, s_70__6_, s_70__5_, s_70__4_, s_70__3_,
         s_70__2_, s_70__1_, s_70__0_, s_71__31_, s_71__30_, s_71__29_,
         s_71__28_, s_71__27_, s_71__26_, s_71__25_, s_71__24_, s_71__23_,
         s_71__22_, s_71__21_, s_71__20_, s_71__19_, s_71__18_, s_71__17_,
         s_71__16_, s_71__15_, s_71__14_, s_71__13_, s_71__12_, s_71__11_,
         s_71__10_, s_71__9_, s_71__8_, s_71__7_, s_71__6_, s_71__5_, s_71__4_,
         s_71__3_, s_71__2_, s_71__1_, s_71__0_, s_72__31_, s_72__30_,
         s_72__29_, s_72__28_, s_72__27_, s_72__26_, s_72__25_, s_72__24_,
         s_72__23_, s_72__22_, s_72__21_, s_72__20_, s_72__19_, s_72__18_,
         s_72__17_, s_72__16_, s_72__15_, s_72__14_, s_72__13_, s_72__12_,
         s_72__11_, s_72__10_, s_72__9_, s_72__8_, s_72__7_, s_72__6_,
         s_72__5_, s_72__4_, s_72__3_, s_72__2_, s_72__1_, s_72__0_, s_73__31_,
         s_73__30_, s_73__29_, s_73__28_, s_73__27_, s_73__26_, s_73__25_,
         s_73__24_, s_73__23_, s_73__22_, s_73__21_, s_73__20_, s_73__19_,
         s_73__18_, s_73__17_, s_73__16_, s_73__15_, s_73__14_, s_73__13_,
         s_73__12_, s_73__11_, s_73__10_, s_73__9_, s_73__8_, s_73__7_,
         s_73__6_, s_73__5_, s_73__4_, s_73__3_, s_73__2_, s_73__1_, s_73__0_,
         s_74__31_, s_74__30_, s_74__29_, s_74__28_, s_74__27_, s_74__26_,
         s_74__25_, s_74__24_, s_74__23_, s_74__22_, s_74__21_, s_74__20_,
         s_74__19_, s_74__18_, s_74__17_, s_74__16_, s_74__15_, s_74__14_,
         s_74__13_, s_74__12_, s_74__11_, s_74__10_, s_74__9_, s_74__8_,
         s_74__7_, s_74__6_, s_74__5_, s_74__4_, s_74__3_, s_74__2_, s_74__1_,
         s_74__0_, s_75__31_, s_75__30_, s_75__29_, s_75__28_, s_75__27_,
         s_75__26_, s_75__25_, s_75__24_, s_75__23_, s_75__22_, s_75__21_,
         s_75__20_, s_75__19_, s_75__18_, s_75__17_, s_75__16_, s_75__15_,
         s_75__14_, s_75__13_, s_75__12_, s_75__11_, s_75__10_, s_75__9_,
         s_75__8_, s_75__7_, s_75__6_, s_75__5_, s_75__4_, s_75__3_, s_75__2_,
         s_75__1_, s_75__0_, s_76__31_, s_76__30_, s_76__29_, s_76__28_,
         s_76__27_, s_76__26_, s_76__25_, s_76__24_, s_76__23_, s_76__22_,
         s_76__21_, s_76__20_, s_76__19_, s_76__18_, s_76__17_, s_76__16_,
         s_76__15_, s_76__14_, s_76__13_, s_76__12_, s_76__11_, s_76__10_,
         s_76__9_, s_76__8_, s_76__7_, s_76__6_, s_76__5_, s_76__4_, s_76__3_,
         s_76__2_, s_76__1_, s_76__0_, s_77__31_, s_77__30_, s_77__29_,
         s_77__28_, s_77__27_, s_77__26_, s_77__25_, s_77__24_, s_77__23_,
         s_77__22_, s_77__21_, s_77__20_, s_77__19_, s_77__18_, s_77__17_,
         s_77__16_, s_77__15_, s_77__14_, s_77__13_, s_77__12_, s_77__11_,
         s_77__10_, s_77__9_, s_77__8_, s_77__7_, s_77__6_, s_77__5_, s_77__4_,
         s_77__3_, s_77__2_, s_77__1_, s_77__0_, s_78__31_, s_78__30_,
         s_78__29_, s_78__28_, s_78__27_, s_78__26_, s_78__25_, s_78__24_,
         s_78__23_, s_78__22_, s_78__21_, s_78__20_, s_78__19_, s_78__18_,
         s_78__17_, s_78__16_, s_78__15_, s_78__14_, s_78__13_, s_78__12_,
         s_78__11_, s_78__10_, s_78__9_, s_78__8_, s_78__7_, s_78__6_,
         s_78__5_, s_78__4_, s_78__3_, s_78__2_, s_78__1_, s_78__0_, s_79__31_,
         s_79__30_, s_79__29_, s_79__28_, s_79__27_, s_79__26_, s_79__25_,
         s_79__24_, s_79__23_, s_79__22_, s_79__21_, s_79__20_, s_79__19_,
         s_79__18_, s_79__17_, s_79__16_, s_79__15_, s_79__14_, s_79__13_,
         s_79__12_, s_79__11_, s_79__10_, s_79__9_, s_79__8_, s_79__7_,
         s_79__6_, s_79__5_, s_79__4_, s_79__3_, s_79__2_, s_79__1_, s_79__0_,
         n1, n2, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32;
  wire   [479:0] sr;

  reg_24 R_0 ( .Reset(n1293), .Clk(Clk), .Load(n2), .Din(Output), .Dout({
        y_1__31_, y_1__30_, y_1__29_, y_1__28_, y_1__27_, y_1__26_, y_1__25_, 
        y_1__24_, y_1__23_, y_1__22_, y_1__21_, y_1__20_, y_1__19_, y_1__18_, 
        y_1__17_, y_1__16_, y_1__15_, y_1__14_, y_1__13_, y_1__12_, y_1__11_, 
        y_1__10_, y_1__9_, y_1__8_, y_1__7_, y_1__6_, y_1__5_, y_1__4_, 
        y_1__3_, y_1__2_, y_1__1_, y_1__0_}) );
  reg_23 R_1 ( .Reset(n1297), .Clk(Clk), .Load(n2), .Din({y_1__31_, y_1__30_, 
        y_1__29_, y_1__28_, y_1__27_, y_1__26_, y_1__25_, y_1__24_, y_1__23_, 
        y_1__22_, n1181, y_1__20_, n1184, n1183, n1198, n1215, n1203, n1214, 
        n1211, n1209, n1222, y_1__10_, n1225, n1218, n1229, n1188, n1228, 
        n1217, n1226, n1220, n1213, n1189}), .Dout({y_2__31_, y_2__30_, 
        y_2__29_, y_2__28_, y_2__27_, y_2__26_, y_2__25_, y_2__24_, y_2__23_, 
        y_2__22_, y_2__21_, y_2__20_, y_2__19_, y_2__18_, y_2__17_, y_2__16_, 
        y_2__15_, y_2__14_, y_2__13_, y_2__12_, y_2__11_, y_2__10_, y_2__9_, 
        y_2__8_, y_2__7_, y_2__6_, y_2__5_, y_2__4_, y_2__3_, y_2__2_, y_2__1_, 
        y_2__0_}) );
  reg_22 R_2 ( .Reset(n1297), .Clk(Clk), .Load(n2), .Din({y_2__31_, y_2__30_, 
        y_2__29_, y_2__28_, y_2__27_, y_2__26_, y_2__25_, y_2__24_, y_2__23_, 
        y_2__22_, n1292, n1289, n1285, n1283, n1281, n1278, n1275, n1272, 
        n1269, n1266, n1263, n1260, n1258, n1255, n1252, n1250, n1247, n1244, 
        n1240, n1238, n1234, n1232}), .Dout({y_3__31_, y_3__30_, y_3__29_, 
        y_3__28_, y_3__27_, y_3__26_, y_3__25_, y_3__24_, y_3__23_, y_3__22_, 
        y_3__21_, y_3__20_, y_3__19_, y_3__18_, y_3__17_, y_3__16_, y_3__15_, 
        y_3__14_, y_3__13_, y_3__12_, y_3__11_, y_3__10_, y_3__9_, y_3__8_, 
        y_3__7_, y_3__6_, y_3__5_, y_3__4_, y_3__3_, y_3__2_, y_3__1_, y_3__0_}) );
  reg_21 R_3 ( .Reset(n1298), .Clk(Clk), .Load(n2), .Din({y_3__31_, y_3__30_, 
        y_3__29_, y_3__28_, y_3__27_, y_3__26_, y_3__25_, y_3__24_, y_3__23_, 
        y_3__22_, y_3__21_, y_3__20_, y_3__19_, y_3__18_, y_3__17_, y_3__16_, 
        y_3__15_, y_3__14_, n1200, y_3__12_, n1187, y_3__10_, y_3__9_, y_3__8_, 
        y_3__7_, y_3__6_, y_3__5_, y_3__4_, y_3__3_, y_3__2_, y_3__1_, y_3__0_}), .Dout({y_4__31_, y_4__30_, y_4__29_, y_4__28_, y_4__27_, y_4__26_, y_4__25_, 
        y_4__24_, y_4__23_, y_4__22_, y_4__21_, y_4__20_, y_4__19_, y_4__18_, 
        y_4__17_, y_4__16_, y_4__15_, y_4__14_, y_4__13_, y_4__12_, y_4__11_, 
        y_4__10_, y_4__9_, y_4__8_, y_4__7_, y_4__6_, y_4__5_, y_4__4_, 
        y_4__3_, y_4__2_, y_4__1_, y_4__0_}) );
  reg_20 R_4 ( .Reset(n1298), .Clk(Clk), .Load(n2), .Din({y_4__31_, y_4__30_, 
        y_4__29_, y_4__28_, y_4__27_, y_4__26_, y_4__25_, y_4__24_, y_4__23_, 
        y_4__22_, y_4__21_, y_4__20_, y_4__19_, y_4__18_, y_4__17_, y_4__16_, 
        y_4__15_, y_4__14_, n1201, y_4__12_, n1196, y_4__10_, y_4__9_, n1180, 
        y_4__7_, y_4__6_, n1194, n1182, y_4__3_, y_4__2_, y_4__1_, y_4__0_}), 
        .Dout({y_5__31_, y_5__30_, y_5__29_, y_5__28_, y_5__27_, y_5__26_, 
        y_5__25_, y_5__24_, y_5__23_, y_5__22_, y_5__21_, y_5__20_, y_5__19_, 
        y_5__18_, y_5__17_, y_5__16_, y_5__15_, y_5__14_, y_5__13_, y_5__12_, 
        y_5__11_, y_5__10_, y_5__9_, y_5__8_, y_5__7_, y_5__6_, y_5__5_, 
        y_5__4_, y_5__3_, y_5__2_, y_5__1_, y_5__0_}) );
  reg_19 R_5 ( .Reset(n1299), .Clk(Clk), .Load(n2), .Din({y_5__31_, y_5__30_, 
        y_5__29_, y_5__28_, y_5__27_, y_5__26_, y_5__25_, y_5__24_, y_5__23_, 
        y_5__22_, y_5__21_, y_5__20_, y_5__19_, y_5__18_, y_5__17_, y_5__16_, 
        y_5__15_, y_5__14_, y_5__13_, y_5__12_, y_5__11_, y_5__10_, n1178, 
        y_5__8_, y_5__7_, y_5__6_, y_5__5_, y_5__4_, y_5__3_, y_5__2_, y_5__1_, 
        y_5__0_}), .Dout({y_6__31_, y_6__30_, y_6__29_, y_6__28_, y_6__27_, 
        y_6__26_, y_6__25_, y_6__24_, y_6__23_, y_6__22_, y_6__21_, y_6__20_, 
        y_6__19_, y_6__18_, y_6__17_, y_6__16_, y_6__15_, y_6__14_, y_6__13_, 
        y_6__12_, y_6__11_, y_6__10_, y_6__9_, y_6__8_, y_6__7_, y_6__6_, 
        y_6__5_, y_6__4_, y_6__3_, y_6__2_, y_6__1_, y_6__0_}) );
  reg_18 R_6 ( .Reset(n1299), .Clk(Clk), .Load(n2), .Din({y_6__31_, y_6__30_, 
        y_6__29_, y_6__28_, y_6__27_, y_6__26_, y_6__25_, y_6__24_, y_6__23_, 
        y_6__22_, y_6__21_, y_6__20_, y_6__19_, y_6__18_, y_6__17_, y_6__16_, 
        y_6__15_, y_6__14_, y_6__13_, y_6__12_, y_6__11_, y_6__10_, y_6__9_, 
        y_6__8_, y_6__7_, y_6__6_, y_6__5_, y_6__4_, y_6__3_, y_6__2_, y_6__1_, 
        y_6__0_}), .Dout({y_7__31_, y_7__30_, y_7__29_, y_7__28_, y_7__27_, 
        y_7__26_, y_7__25_, y_7__24_, y_7__23_, y_7__22_, y_7__21_, y_7__20_, 
        y_7__19_, y_7__18_, y_7__17_, y_7__16_, y_7__15_, y_7__14_, y_7__13_, 
        y_7__12_, y_7__11_, y_7__10_, y_7__9_, y_7__8_, y_7__7_, y_7__6_, 
        y_7__5_, y_7__4_, y_7__3_, y_7__2_, y_7__1_, y_7__0_}) );
  reg_17 R_7 ( .Reset(n1299), .Clk(Clk), .Load(n2), .Din({y_7__31_, y_7__30_, 
        y_7__29_, y_7__28_, y_7__27_, y_7__26_, y_7__25_, y_7__24_, y_7__23_, 
        y_7__22_, y_7__21_, y_7__20_, y_7__19_, y_7__18_, y_7__17_, y_7__16_, 
        y_7__15_, y_7__14_, y_7__13_, y_7__12_, y_7__11_, y_7__10_, y_7__9_, 
        y_7__8_, y_7__7_, y_7__6_, y_7__5_, y_7__4_, y_7__3_, y_7__2_, y_7__1_, 
        y_7__0_}), .Dout({y_8__31_, y_8__30_, y_8__29_, y_8__28_, y_8__27_, 
        y_8__26_, y_8__25_, y_8__24_, y_8__23_, y_8__22_, y_8__21_, y_8__20_, 
        y_8__19_, y_8__18_, y_8__17_, y_8__16_, y_8__15_, y_8__14_, y_8__13_, 
        y_8__12_, y_8__11_, y_8__10_, y_8__9_, y_8__8_, y_8__7_, y_8__6_, 
        y_8__5_, y_8__4_, y_8__3_, y_8__2_, y_8__1_, y_8__0_}) );
  reg_16 R_8 ( .Reset(n1298), .Clk(Clk), .Load(n2), .Din({y_8__31_, y_8__30_, 
        y_8__29_, y_8__28_, y_8__27_, y_8__26_, y_8__25_, y_8__24_, y_8__23_, 
        y_8__22_, y_8__21_, y_8__20_, y_8__19_, y_8__18_, y_8__17_, y_8__16_, 
        y_8__15_, y_8__14_, y_8__13_, y_8__12_, y_8__11_, y_8__10_, y_8__9_, 
        y_8__8_, y_8__7_, y_8__6_, y_8__5_, y_8__4_, y_8__3_, y_8__2_, y_8__1_, 
        y_8__0_}), .Dout({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32}) );
  adder_0 S92 ( .A({s_91__31_, s_91__30_, s_91__29_, s_91__28_, s_91__27_, 
        s_91__26_, s_91__25_, s_91__24_, s_91__23_, s_91__22_, s_91__21_, 
        s_91__20_, s_91__19_, s_91__18_, s_91__17_, s_91__16_, s_91__15_, 
        s_91__14_, s_91__13_, s_91__12_, s_91__11_, s_91__10_, s_91__9_, 
        s_91__8_, s_91__7_, s_91__6_, s_91__5_, s_91__4_, s_91__3_, s_91__2_, 
        s_91__1_, s_91__0_}), .B({s_90__31_, s_90__30_, s_90__29_, s_90__28_, 
        s_90__27_, s_90__26_, s_90__25_, s_90__24_, s_90__23_, s_90__22_, 
        s_90__21_, s_90__20_, s_90__19_, s_90__18_, s_90__17_, s_90__16_, 
        s_90__15_, s_90__14_, s_90__13_, s_90__12_, s_90__11_, s_90__10_, 
        s_90__9_, s_90__8_, s_90__7_, s_90__6_, s_90__5_, s_90__4_, s_90__3_, 
        s_90__2_, s_90__1_, s_90__0_}), .O(Output) );
  reg_15 R0 ( .Reset(n1297), .Clk(Clk), .Load(n2), .Din({s_89__31_, s_89__30_, 
        s_89__29_, s_89__28_, s_89__27_, s_89__26_, s_89__25_, s_89__24_, 
        s_89__23_, s_89__22_, s_89__21_, s_89__20_, s_89__19_, s_89__18_, 
        s_89__17_, s_89__16_, s_89__15_, s_89__14_, s_89__13_, s_89__12_, 
        s_89__11_, s_89__10_, s_89__9_, s_89__8_, s_89__7_, s_89__6_, s_89__5_, 
        s_89__4_, s_89__3_, s_89__2_, s_89__1_, s_89__0_}), .Dout(sr[479:448])
         );
  reg_14 R1 ( .Reset(n1295), .Clk(Clk), .Load(n2), .Din({s_88__31_, s_88__30_, 
        s_88__29_, s_88__28_, s_88__27_, s_88__26_, s_88__25_, s_88__24_, 
        s_88__23_, s_88__22_, s_88__21_, s_88__20_, s_88__19_, s_88__18_, 
        s_88__17_, s_88__16_, s_88__15_, s_88__14_, s_88__13_, s_88__12_, 
        s_88__11_, s_88__10_, s_88__9_, s_88__8_, s_88__7_, s_88__6_, s_88__5_, 
        s_88__4_, s_88__3_, s_88__2_, s_88__1_, s_88__0_}), .Dout(sr[447:416])
         );
  adder_45 S91 ( .A(sr[479:448]), .B(sr[447:416]), .O({s_91__31_, s_91__30_, 
        s_91__29_, s_91__28_, s_91__27_, s_91__26_, s_91__25_, s_91__24_, 
        s_91__23_, s_91__22_, s_91__21_, s_91__20_, s_91__19_, s_91__18_, 
        s_91__17_, s_91__16_, s_91__15_, s_91__14_, s_91__13_, s_91__12_, 
        s_91__11_, s_91__10_, s_91__9_, s_91__8_, s_91__7_, s_91__6_, s_91__5_, 
        s_91__4_, s_91__3_, s_91__2_, s_91__1_, s_91__0_}) );
  adder_44 S89 ( .A({s_85__31_, s_85__30_, s_85__29_, s_85__28_, s_85__27_, 
        s_85__26_, s_85__25_, s_85__24_, s_85__23_, s_85__22_, s_85__21_, 
        s_85__20_, s_85__19_, s_85__18_, s_85__17_, s_85__16_, s_85__15_, 
        s_85__14_, s_85__13_, s_85__12_, s_85__11_, s_85__10_, s_85__9_, 
        s_85__8_, s_85__7_, s_85__6_, s_85__5_, s_85__4_, s_85__3_, s_85__2_, 
        s_85__1_, s_85__0_}), .B({s_84__31_, s_84__30_, s_84__29_, s_84__28_, 
        s_84__27_, s_84__26_, s_84__25_, s_84__24_, s_84__23_, s_84__22_, 
        s_84__21_, s_84__20_, s_84__19_, s_84__18_, s_84__17_, s_84__16_, 
        s_84__15_, s_84__14_, s_84__13_, s_84__12_, s_84__11_, s_84__10_, 
        s_84__9_, s_84__8_, s_84__7_, s_84__6_, s_84__5_, s_84__4_, s_84__3_, 
        s_84__2_, s_84__1_, s_84__0_}), .O({s_89__31_, s_89__30_, s_89__29_, 
        s_89__28_, s_89__27_, s_89__26_, s_89__25_, s_89__24_, s_89__23_, 
        s_89__22_, s_89__21_, s_89__20_, s_89__19_, s_89__18_, s_89__17_, 
        s_89__16_, s_89__15_, s_89__14_, s_89__13_, s_89__12_, s_89__11_, 
        s_89__10_, s_89__9_, s_89__8_, s_89__7_, s_89__6_, s_89__5_, s_89__4_, 
        s_89__3_, s_89__2_, s_89__1_, s_89__0_}) );
  adder_43 S85 ( .A({y_2__25_, y_2__24_, y_2__23_, y_2__22_, n1292, n1289, 
        n1286, n1283, n1281, n1279, n1276, n1273, n1270, n1267, n1264, n1261, 
        n1258, n1255, n1253, n1250, n1247, n1244, n1241, n1238, n1234, n1231, 
        n1, n1, n1, n1, n1, n1}), .B({y_1__27_, y_1__26_, y_1__25_, y_1__24_, 
        y_1__23_, y_1__22_, n1181, y_1__20_, n1184, n1183, n1198, n1215, n1203, 
        n1214, n1211, n1209, n1222, y_1__10_, n1225, n1218, n1229, n1188, 
        n1228, n1217, n1226, n1220, n1213, y_1__0_, n1, n1, n1, n1}), .O({
        s_85__31_, s_85__30_, s_85__29_, s_85__28_, s_85__27_, s_85__26_, 
        s_85__25_, s_85__24_, s_85__23_, s_85__22_, s_85__21_, s_85__20_, 
        s_85__19_, s_85__18_, s_85__17_, s_85__16_, s_85__15_, s_85__14_, 
        s_85__13_, s_85__12_, s_85__11_, s_85__10_, s_85__9_, s_85__8_, 
        s_85__7_, s_85__6_, s_85__5_, s_85__4_, s_85__3_, s_85__2_, s_85__1_, 
        s_85__0_}) );
  adder_42 S84 ( .A({y_2__29_, y_2__28_, y_2__27_, y_2__26_, y_2__25_, 
        y_2__24_, y_2__23_, y_2__22_, n1292, n1289, n1285, n1283, n1281, n1278, 
        n1275, n1272, n1269, n1266, n1263, n1260, n1257, n1255, n1252, n1250, 
        n1247, n1244, n1240, n1238, n1235, n1232, n1, n1}), .B({y_2__28_, 
        y_2__27_, y_2__26_, y_2__25_, y_2__24_, y_2__23_, y_2__22_, n1291, 
        n1288, n1286, n1283, n1281, n1278, n1276, n1272, n1270, n1267, n1263, 
        n1260, n1258, n1255, n1253, n1249, n1246, n1243, n1240, n1237, n1235, 
        n1231, n1, n1, n1}), .O({s_84__31_, s_84__30_, s_84__29_, s_84__28_, 
        s_84__27_, s_84__26_, s_84__25_, s_84__24_, s_84__23_, s_84__22_, 
        s_84__21_, s_84__20_, s_84__19_, s_84__18_, s_84__17_, s_84__16_, 
        s_84__15_, s_84__14_, s_84__13_, s_84__12_, s_84__11_, s_84__10_, 
        s_84__9_, s_84__8_, s_84__7_, s_84__6_, s_84__5_, s_84__4_, s_84__3_, 
        s_84__2_, s_84__1_, s_84__0_}) );
  adder_41 S88 ( .A({s_87__31_, s_87__30_, s_87__29_, s_87__28_, s_87__27_, 
        s_87__26_, s_87__25_, s_87__24_, s_87__23_, s_87__22_, s_87__21_, 
        s_87__20_, s_87__19_, s_87__18_, s_87__17_, s_87__16_, s_87__15_, 
        s_87__14_, s_87__13_, s_87__12_, s_87__11_, s_87__10_, s_87__9_, 
        s_87__8_, s_87__7_, s_87__6_, s_87__5_, s_87__4_, s_87__3_, s_87__2_, 
        s_87__1_, s_87__0_}), .B({s_86__31_, s_86__30_, s_86__29_, s_86__28_, 
        s_86__27_, s_86__26_, s_86__25_, s_86__24_, s_86__23_, s_86__22_, 
        s_86__21_, s_86__20_, s_86__19_, s_86__18_, s_86__17_, s_86__16_, 
        s_86__15_, s_86__14_, s_86__13_, s_86__12_, s_86__11_, s_86__10_, 
        s_86__9_, s_86__8_, s_86__7_, s_86__6_, s_86__5_, s_86__4_, s_86__3_, 
        s_86__2_, s_86__1_, s_86__0_}), .O({s_88__31_, s_88__30_, s_88__29_, 
        s_88__28_, s_88__27_, s_88__26_, s_88__25_, s_88__24_, s_88__23_, 
        s_88__22_, s_88__21_, s_88__20_, s_88__19_, s_88__18_, s_88__17_, 
        s_88__16_, s_88__15_, s_88__14_, s_88__13_, s_88__12_, s_88__11_, 
        s_88__10_, s_88__9_, s_88__8_, s_88__7_, s_88__6_, s_88__5_, s_88__4_, 
        s_88__3_, s_88__2_, s_88__1_, s_88__0_}) );
  reg_13 R2 ( .Reset(n1294), .Clk(Clk), .Load(n2), .Din({s_82__31_, s_82__30_, 
        s_82__29_, s_82__28_, s_82__27_, s_82__26_, s_82__25_, s_82__24_, 
        s_82__23_, s_82__22_, s_82__21_, s_82__20_, s_82__19_, s_82__18_, 
        s_82__17_, s_82__16_, s_82__15_, s_82__14_, s_82__13_, s_82__12_, 
        s_82__11_, s_82__10_, s_82__9_, s_82__8_, s_82__7_, s_82__6_, s_82__5_, 
        s_82__4_, s_82__3_, s_82__2_, s_82__1_, s_82__0_}), .Dout(sr[415:384])
         );
  reg_12 R3 ( .Reset(n1295), .Clk(Clk), .Load(n2), .Din({s_81__31_, s_81__30_, 
        s_81__29_, s_81__28_, s_81__27_, s_81__26_, s_81__25_, s_81__24_, 
        s_81__23_, s_81__22_, s_81__21_, s_81__20_, s_81__19_, s_81__18_, 
        s_81__17_, s_81__16_, s_81__15_, s_81__14_, s_81__13_, s_81__12_, 
        s_81__11_, s_81__10_, s_81__9_, s_81__8_, s_81__7_, s_81__6_, s_81__5_, 
        s_81__4_, s_81__3_, s_81__2_, s_81__1_, s_81__0_}), .Dout(sr[383:352])
         );
  adder_40 S87 ( .A(sr[415:384]), .B(sr[383:352]), .O({s_87__31_, s_87__30_, 
        s_87__29_, s_87__28_, s_87__27_, s_87__26_, s_87__25_, s_87__24_, 
        s_87__23_, s_87__22_, s_87__21_, s_87__20_, s_87__19_, s_87__18_, 
        s_87__17_, s_87__16_, s_87__15_, s_87__14_, s_87__13_, s_87__12_, 
        s_87__11_, s_87__10_, s_87__9_, s_87__8_, s_87__7_, s_87__6_, s_87__5_, 
        s_87__4_, s_87__3_, s_87__2_, s_87__1_, s_87__0_}) );
  adder_39 S82 ( .A({s_78__31_, s_78__30_, s_78__29_, s_78__28_, s_78__27_, 
        s_78__26_, s_78__25_, s_78__24_, s_78__23_, s_78__22_, s_78__21_, 
        s_78__20_, s_78__19_, s_78__18_, s_78__17_, s_78__16_, s_78__15_, 
        s_78__14_, s_78__13_, s_78__12_, s_78__11_, s_78__10_, s_78__9_, 
        s_78__8_, s_78__7_, s_78__6_, s_78__5_, s_78__4_, s_78__3_, s_78__2_, 
        s_78__1_, s_78__0_}), .B({s_77__31_, s_77__30_, s_77__29_, s_77__28_, 
        s_77__27_, s_77__26_, s_77__25_, s_77__24_, s_77__23_, s_77__22_, 
        s_77__21_, s_77__20_, s_77__19_, s_77__18_, s_77__17_, s_77__16_, 
        s_77__15_, s_77__14_, s_77__13_, s_77__12_, s_77__11_, s_77__10_, 
        s_77__9_, s_77__8_, s_77__7_, s_77__6_, s_77__5_, s_77__4_, s_77__3_, 
        s_77__2_, s_77__1_, s_77__0_}), .O({s_82__31_, s_82__30_, s_82__29_, 
        s_82__28_, s_82__27_, s_82__26_, s_82__25_, s_82__24_, s_82__23_, 
        s_82__22_, s_82__21_, s_82__20_, s_82__19_, s_82__18_, s_82__17_, 
        s_82__16_, s_82__15_, s_82__14_, s_82__13_, s_82__12_, s_82__11_, 
        s_82__10_, s_82__9_, s_82__8_, s_82__7_, s_82__6_, s_82__5_, s_82__4_, 
        s_82__3_, s_82__2_, s_82__1_, s_82__0_}) );
  reg_11 R4 ( .Reset(n1294), .Clk(Clk), .Load(n2), .Din({s_71__31_, s_71__30_, 
        s_71__29_, s_71__28_, s_71__27_, s_71__26_, s_71__25_, s_71__24_, 
        s_71__23_, s_71__22_, s_71__21_, s_71__20_, s_71__19_, s_71__18_, 
        s_71__17_, s_71__16_, s_71__15_, s_71__14_, s_71__13_, s_71__12_, 
        s_71__11_, s_71__10_, s_71__9_, s_71__8_, s_71__7_, s_71__6_, s_71__5_, 
        s_71__4_, s_71__3_, s_71__2_, s_71__1_, s_71__0_}), .Dout(sr[351:320])
         );
  reg_10 R5 ( .Reset(n1299), .Clk(Clk), .Load(n2), .Din({s_70__31_, s_70__30_, 
        s_70__29_, s_70__28_, s_70__27_, s_70__26_, s_70__25_, s_70__24_, 
        s_70__23_, s_70__22_, s_70__21_, s_70__20_, s_70__19_, s_70__18_, 
        s_70__17_, s_70__16_, s_70__15_, s_70__14_, s_70__13_, s_70__12_, 
        s_70__11_, s_70__10_, s_70__9_, s_70__8_, s_70__7_, s_70__6_, s_70__5_, 
        s_70__4_, s_70__3_, s_70__2_, s_70__1_, s_70__0_}), .Dout(sr[319:288])
         );
  adder_38 S78 ( .A(sr[351:320]), .B(sr[319:288]), .O({s_78__31_, s_78__30_, 
        s_78__29_, s_78__28_, s_78__27_, s_78__26_, s_78__25_, s_78__24_, 
        s_78__23_, s_78__22_, s_78__21_, s_78__20_, s_78__19_, s_78__18_, 
        s_78__17_, s_78__16_, s_78__15_, s_78__14_, s_78__13_, s_78__12_, 
        s_78__11_, s_78__10_, s_78__9_, s_78__8_, s_78__7_, s_78__6_, s_78__5_, 
        s_78__4_, s_78__3_, s_78__2_, s_78__1_, s_78__0_}) );
  adder_37 S71 ( .A({s_55__31_, s_55__30_, s_55__29_, s_55__28_, s_55__27_, 
        s_55__26_, s_55__25_, s_55__24_, s_55__23_, s_55__22_, s_55__21_, 
        s_55__20_, s_55__19_, s_55__18_, s_55__17_, s_55__16_, s_55__15_, 
        s_55__14_, s_55__13_, s_55__12_, s_55__11_, s_55__10_, s_55__9_, 
        s_55__8_, s_55__7_, s_55__6_, s_55__5_, s_55__4_, s_55__3_, s_55__2_, 
        s_55__1_, s_55__0_}), .B({s_54__31_, s_54__30_, s_54__29_, s_54__28_, 
        s_54__27_, s_54__26_, s_54__25_, s_54__24_, s_54__23_, s_54__22_, 
        s_54__21_, s_54__20_, s_54__19_, s_54__18_, s_54__17_, s_54__16_, 
        s_54__15_, s_54__14_, s_54__13_, s_54__12_, s_54__11_, s_54__10_, 
        s_54__9_, s_54__8_, s_54__7_, s_54__6_, s_54__5_, s_54__4_, s_54__3_, 
        s_54__2_, s_54__1_, s_54__0_}), .O({s_71__31_, s_71__30_, s_71__29_, 
        s_71__28_, s_71__27_, s_71__26_, s_71__25_, s_71__24_, s_71__23_, 
        s_71__22_, s_71__21_, s_71__20_, s_71__19_, s_71__18_, s_71__17_, 
        s_71__16_, s_71__15_, s_71__14_, s_71__13_, s_71__12_, s_71__11_, 
        s_71__10_, s_71__9_, s_71__8_, s_71__7_, s_71__6_, s_71__5_, s_71__4_, 
        s_71__3_, s_71__2_, s_71__1_, s_71__0_}) );
  adder_36 S55 ( .A({Input[180:160], n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1}), .B({y_5__27_, y_5__26_, y_5__25_, y_5__24_, y_5__23_, y_5__22_, 
        y_5__21_, y_5__20_, y_5__19_, y_5__18_, y_5__17_, y_5__16_, y_5__15_, 
        y_5__14_, y_5__13_, y_5__12_, y_5__11_, y_5__10_, n1178, y_5__8_, 
        y_5__7_, y_5__6_, y_5__5_, y_5__4_, y_5__3_, y_5__2_, y_5__1_, y_5__0_, 
        n1, n1, n1, n1}), .O({s_55__31_, s_55__30_, s_55__29_, s_55__28_, 
        s_55__27_, s_55__26_, s_55__25_, s_55__24_, s_55__23_, s_55__22_, 
        s_55__21_, s_55__20_, s_55__19_, s_55__18_, s_55__17_, s_55__16_, 
        s_55__15_, s_55__14_, s_55__13_, s_55__12_, s_55__11_, s_55__10_, 
        s_55__9_, s_55__8_, s_55__7_, s_55__6_, s_55__5_, s_55__4_, s_55__3_, 
        s_55__2_, s_55__1_, s_55__0_}) );
  adder_35 S54 ( .A(Input[191:160]), .B({Input[181:160], n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1}), .O({s_54__31_, s_54__30_, s_54__29_, s_54__28_, 
        s_54__27_, s_54__26_, s_54__25_, s_54__24_, s_54__23_, s_54__22_, 
        s_54__21_, s_54__20_, s_54__19_, s_54__18_, s_54__17_, s_54__16_, 
        s_54__15_, s_54__14_, s_54__13_, s_54__12_, s_54__11_, s_54__10_, 
        s_54__9_, s_54__8_, s_54__7_, s_54__6_, s_54__5_, s_54__4_, s_54__3_, 
        s_54__2_, s_54__1_, s_54__0_}) );
  adder_34 S70 ( .A({s_57__31_, s_57__30_, s_57__29_, s_57__28_, s_57__27_, 
        s_57__26_, s_57__25_, s_57__24_, s_57__23_, s_57__22_, s_57__21_, 
        s_57__20_, s_57__19_, s_57__18_, s_57__17_, s_57__16_, s_57__15_, 
        s_57__14_, s_57__13_, s_57__12_, s_57__11_, s_57__10_, s_57__9_, 
        s_57__8_, s_57__7_, s_57__6_, s_57__5_, s_57__4_, s_57__3_, s_57__2_, 
        s_57__1_, s_57__0_}), .B({s_56__31_, s_56__30_, s_56__29_, s_56__28_, 
        s_56__27_, s_56__26_, s_56__25_, s_56__24_, s_56__23_, s_56__22_, 
        s_56__21_, s_56__20_, s_56__19_, s_56__18_, s_56__17_, s_56__16_, 
        s_56__15_, s_56__14_, s_56__13_, s_56__12_, s_56__11_, s_56__10_, 
        s_56__9_, s_56__8_, s_56__7_, s_56__6_, s_56__5_, s_56__4_, s_56__3_, 
        s_56__2_, s_56__1_, s_56__0_}), .O({s_70__31_, s_70__30_, s_70__29_, 
        s_70__28_, s_70__27_, s_70__26_, s_70__25_, s_70__24_, s_70__23_, 
        s_70__22_, s_70__21_, s_70__20_, s_70__19_, s_70__18_, s_70__17_, 
        s_70__16_, s_70__15_, s_70__14_, s_70__13_, s_70__12_, s_70__11_, 
        s_70__10_, s_70__9_, s_70__8_, s_70__7_, s_70__6_, s_70__5_, s_70__4_, 
        s_70__3_, s_70__2_, s_70__1_, s_70__0_}) );
  adder_33 S57 ( .A({Input[215:192], n1, n1, n1, n1, n1, n1, n1, n1}), .B({
        y_4__29_, y_4__28_, y_4__27_, y_4__26_, y_4__25_, y_4__24_, y_4__23_, 
        y_4__22_, y_4__21_, y_4__20_, y_4__19_, y_4__18_, y_4__17_, y_4__16_, 
        y_4__15_, y_4__14_, y_4__13_, y_4__12_, n1196, y_4__10_, y_4__9_, 
        n1180, y_4__7_, y_4__6_, y_4__5_, n1182, y_4__3_, y_4__2_, y_4__1_, 
        y_4__0_, n1, n1}), .O({s_57__31_, s_57__30_, s_57__29_, s_57__28_, 
        s_57__27_, s_57__26_, s_57__25_, s_57__24_, s_57__23_, s_57__22_, 
        s_57__21_, s_57__20_, s_57__19_, s_57__18_, s_57__17_, s_57__16_, 
        s_57__15_, s_57__14_, s_57__13_, s_57__12_, s_57__11_, s_57__10_, 
        s_57__9_, s_57__8_, s_57__7_, s_57__6_, s_57__5_, s_57__4_, s_57__3_, 
        s_57__2_, s_57__1_, s_57__0_}) );
  adder_32 S56 ( .A({y_5__26_, y_5__25_, y_5__24_, y_5__23_, y_5__22_, 
        y_5__21_, y_5__20_, y_5__19_, y_5__18_, y_5__17_, y_5__16_, y_5__15_, 
        y_5__14_, y_5__13_, y_5__12_, y_5__11_, y_5__10_, n1178, y_5__8_, 
        y_5__7_, y_5__6_, y_5__5_, y_5__4_, y_5__3_, y_5__2_, y_5__1_, y_5__0_, 
        n1, n1, n1, n1, n1}), .B({Input[216:192], n1, n1, n1, n1, n1, n1, n1}), 
        .O({s_56__31_, s_56__30_, s_56__29_, s_56__28_, s_56__27_, s_56__26_, 
        s_56__25_, s_56__24_, s_56__23_, s_56__22_, s_56__21_, s_56__20_, 
        s_56__19_, s_56__18_, s_56__17_, s_56__16_, s_56__15_, s_56__14_, 
        s_56__13_, s_56__12_, s_56__11_, s_56__10_, s_56__9_, s_56__8_, 
        s_56__7_, s_56__6_, s_56__5_, s_56__4_, s_56__3_, s_56__2_, s_56__1_, 
        s_56__0_}) );
  reg_9 R6 ( .Reset(n1295), .Clk(Clk), .Load(n2), .Din({s_73__31_, s_73__30_, 
        s_73__29_, s_73__28_, s_73__27_, s_73__26_, s_73__25_, s_73__24_, 
        s_73__23_, s_73__22_, s_73__21_, s_73__20_, s_73__19_, s_73__18_, 
        s_73__17_, s_73__16_, s_73__15_, s_73__14_, s_73__13_, s_73__12_, 
        s_73__11_, s_73__10_, s_73__9_, s_73__8_, s_73__7_, s_73__6_, s_73__5_, 
        s_73__4_, s_73__3_, s_73__2_, s_73__1_, s_73__0_}), .Dout(sr[287:256])
         );
  reg_8 R7 ( .Reset(n1294), .Clk(Clk), .Load(n2), .Din({s_72__31_, s_72__30_, 
        s_72__29_, s_72__28_, s_72__27_, s_72__26_, s_72__25_, s_72__24_, 
        s_72__23_, s_72__22_, s_72__21_, s_72__20_, s_72__19_, s_72__18_, 
        s_72__17_, s_72__16_, s_72__15_, s_72__14_, s_72__13_, s_72__12_, 
        s_72__11_, s_72__10_, s_72__9_, s_72__8_, s_72__7_, s_72__6_, s_72__5_, 
        s_72__4_, s_72__3_, s_72__2_, s_72__1_, s_72__0_}), .Dout(sr[255:224])
         );
  adder_31 S77 ( .A(sr[287:256]), .B(sr[255:224]), .O({s_77__31_, s_77__30_, 
        s_77__29_, s_77__28_, s_77__27_, s_77__26_, s_77__25_, s_77__24_, 
        s_77__23_, s_77__22_, s_77__21_, s_77__20_, s_77__19_, s_77__18_, 
        s_77__17_, s_77__16_, s_77__15_, s_77__14_, s_77__13_, s_77__12_, 
        s_77__11_, s_77__10_, s_77__9_, s_77__8_, s_77__7_, s_77__6_, s_77__5_, 
        s_77__4_, s_77__3_, s_77__2_, s_77__1_, s_77__0_}) );
  adder_30 S73 ( .A({s_51__31_, s_51__30_, s_51__29_, s_51__28_, s_51__27_, 
        s_51__26_, s_51__25_, s_51__24_, s_51__23_, s_51__22_, s_51__21_, 
        s_51__20_, s_51__19_, s_51__18_, s_51__17_, s_51__16_, s_51__15_, 
        s_51__14_, s_51__13_, s_51__12_, s_51__11_, s_51__10_, s_51__9_, 
        s_51__8_, s_51__7_, s_51__6_, s_51__5_, s_51__4_, s_51__3_, s_51__2_, 
        s_51__1_, s_51__0_}), .B({s_50__31_, s_50__30_, s_50__29_, s_50__28_, 
        s_50__27_, s_50__26_, s_50__25_, s_50__24_, s_50__23_, s_50__22_, 
        s_50__21_, s_50__20_, s_50__19_, s_50__18_, s_50__17_, s_50__16_, 
        s_50__15_, s_50__14_, s_50__13_, s_50__12_, s_50__11_, s_50__10_, 
        s_50__9_, s_50__8_, s_50__7_, s_50__6_, s_50__5_, s_50__4_, s_50__3_, 
        s_50__2_, s_50__1_, s_50__0_}), .O({s_73__31_, s_73__30_, s_73__29_, 
        s_73__28_, s_73__27_, s_73__26_, s_73__25_, s_73__24_, s_73__23_, 
        s_73__22_, s_73__21_, s_73__20_, s_73__19_, s_73__18_, s_73__17_, 
        s_73__16_, s_73__15_, s_73__14_, s_73__13_, s_73__12_, s_73__11_, 
        s_73__10_, s_73__9_, s_73__8_, s_73__7_, s_73__6_, s_73__5_, s_73__4_, 
        s_73__3_, s_73__2_, s_73__1_, s_73__0_}) );
  adder_29 S51 ( .A({Input[119:96], n1, n1, n1, n1, n1, n1, n1, n1}), .B(
        Input[159:128]), .O({s_51__31_, s_51__30_, s_51__29_, s_51__28_, 
        s_51__27_, s_51__26_, s_51__25_, s_51__24_, s_51__23_, s_51__22_, 
        s_51__21_, s_51__20_, s_51__19_, s_51__18_, s_51__17_, s_51__16_, 
        s_51__15_, s_51__14_, s_51__13_, s_51__12_, s_51__11_, s_51__10_, 
        s_51__9_, s_51__8_, s_51__7_, s_51__6_, s_51__5_, s_51__4_, s_51__3_, 
        s_51__2_, s_51__1_, s_51__0_}) );
  adder_28 S50 ( .A({Input[89:68], n1193, Input[66:64], n1, n1, n1, n1, n1, n1}), .B({Input[120:96], n1, n1, n1, n1, n1, n1, n1}), .O({s_50__31_, s_50__30_, 
        s_50__29_, s_50__28_, s_50__27_, s_50__26_, s_50__25_, s_50__24_, 
        s_50__23_, s_50__22_, s_50__21_, s_50__20_, s_50__19_, s_50__18_, 
        s_50__17_, s_50__16_, s_50__15_, s_50__14_, s_50__13_, s_50__12_, 
        s_50__11_, s_50__10_, s_50__9_, s_50__8_, s_50__7_, s_50__6_, s_50__5_, 
        s_50__4_, s_50__3_, s_50__2_, s_50__1_, s_50__0_}) );
  adder_27 S72 ( .A({s_53__31_, s_53__30_, s_53__29_, s_53__28_, s_53__27_, 
        s_53__26_, s_53__25_, s_53__24_, s_53__23_, s_53__22_, s_53__21_, 
        s_53__20_, s_53__19_, s_53__18_, s_53__17_, s_53__16_, s_53__15_, 
        s_53__14_, s_53__13_, s_53__12_, s_53__11_, s_53__10_, s_53__9_, 
        s_53__8_, s_53__7_, s_53__6_, s_53__5_, s_53__4_, s_53__3_, s_53__2_, 
        s_53__1_, s_53__0_}), .B({s_52__31_, s_52__30_, s_52__29_, s_52__28_, 
        s_52__27_, s_52__26_, s_52__25_, s_52__24_, s_52__23_, s_52__22_, 
        s_52__21_, s_52__20_, s_52__19_, s_52__18_, s_52__17_, s_52__16_, 
        s_52__15_, s_52__14_, s_52__13_, s_52__12_, s_52__11_, s_52__10_, 
        s_52__9_, s_52__8_, s_52__7_, s_52__6_, s_52__5_, s_52__4_, s_52__3_, 
        s_52__2_, s_52__1_, s_52__0_}), .O({s_72__31_, s_72__30_, s_72__29_, 
        s_72__28_, s_72__27_, s_72__26_, s_72__25_, s_72__24_, s_72__23_, 
        s_72__22_, s_72__21_, s_72__20_, s_72__19_, s_72__18_, s_72__17_, 
        s_72__16_, s_72__15_, s_72__14_, s_72__13_, s_72__12_, s_72__11_, 
        s_72__10_, s_72__9_, s_72__8_, s_72__7_, s_72__6_, s_72__5_, s_72__4_, 
        s_72__3_, s_72__2_, s_72__1_, s_72__0_}) );
  adder_26 S53 ( .A({y_6__31_, y_6__30_, y_6__29_, y_6__28_, y_6__27_, 
        y_6__26_, y_6__25_, y_6__24_, y_6__23_, y_6__22_, y_6__21_, y_6__20_, 
        y_6__19_, y_6__18_, y_6__17_, y_6__16_, y_6__15_, y_6__14_, y_6__13_, 
        y_6__12_, y_6__11_, y_6__10_, y_6__9_, y_6__8_, y_6__7_, y_6__6_, 
        y_6__5_, y_6__4_, y_6__3_, y_6__2_, y_6__1_, y_6__0_}), .B({y_6__29_, 
        y_6__28_, y_6__27_, y_6__26_, y_6__25_, y_6__24_, y_6__23_, y_6__22_, 
        y_6__21_, y_6__20_, y_6__19_, y_6__18_, y_6__17_, y_6__16_, y_6__15_, 
        y_6__14_, y_6__13_, y_6__12_, y_6__11_, y_6__10_, y_6__9_, y_6__8_, 
        y_6__7_, y_6__6_, y_6__5_, y_6__4_, y_6__3_, y_6__2_, y_6__1_, y_6__0_, 
        n1, n1}), .O({s_53__31_, s_53__30_, s_53__29_, s_53__28_, s_53__27_, 
        s_53__26_, s_53__25_, s_53__24_, s_53__23_, s_53__22_, s_53__21_, 
        s_53__20_, s_53__19_, s_53__18_, s_53__17_, s_53__16_, s_53__15_, 
        s_53__14_, s_53__13_, s_53__12_, s_53__11_, s_53__10_, s_53__9_, 
        s_53__8_, s_53__7_, s_53__6_, s_53__5_, s_53__4_, s_53__3_, s_53__2_, 
        s_53__1_, s_53__0_}) );
  adder_25 S52 ( .A({Input[149:128], n1, n1, n1, n1, n1, n1, n1, n1, n1, n1}), 
        .B({Input[148:128], n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1}), .O({
        s_52__31_, s_52__30_, s_52__29_, s_52__28_, s_52__27_, s_52__26_, 
        s_52__25_, s_52__24_, s_52__23_, s_52__22_, s_52__21_, s_52__20_, 
        s_52__19_, s_52__18_, s_52__17_, s_52__16_, s_52__15_, s_52__14_, 
        s_52__13_, s_52__12_, s_52__11_, s_52__10_, s_52__9_, s_52__8_, 
        s_52__7_, s_52__6_, s_52__5_, s_52__4_, s_52__3_, s_52__2_, s_52__1_, 
        s_52__0_}) );
  adder_24 S81 ( .A({s_80__31_, s_80__30_, s_80__29_, s_80__28_, s_80__27_, 
        s_80__26_, s_80__25_, s_80__24_, s_80__23_, s_80__22_, s_80__21_, 
        s_80__20_, s_80__19_, s_80__18_, s_80__17_, s_80__16_, s_80__15_, 
        s_80__14_, s_80__13_, s_80__12_, s_80__11_, s_80__10_, s_80__9_, 
        s_80__8_, s_80__7_, s_80__6_, s_80__5_, s_80__4_, s_80__3_, s_80__2_, 
        s_80__1_, s_80__0_}), .B({s_79__31_, s_79__30_, s_79__29_, s_79__28_, 
        s_79__27_, s_79__26_, s_79__25_, s_79__24_, s_79__23_, s_79__22_, 
        s_79__21_, s_79__20_, s_79__19_, s_79__18_, s_79__17_, s_79__16_, 
        s_79__15_, s_79__14_, s_79__13_, s_79__12_, s_79__11_, s_79__10_, 
        s_79__9_, s_79__8_, s_79__7_, s_79__6_, s_79__5_, s_79__4_, s_79__3_, 
        s_79__2_, s_79__1_, s_79__0_}), .O({s_81__31_, s_81__30_, s_81__29_, 
        s_81__28_, s_81__27_, s_81__26_, s_81__25_, s_81__24_, s_81__23_, 
        s_81__22_, s_81__21_, s_81__20_, s_81__19_, s_81__18_, s_81__17_, 
        s_81__16_, s_81__15_, s_81__14_, s_81__13_, s_81__12_, s_81__11_, 
        s_81__10_, s_81__9_, s_81__8_, s_81__7_, s_81__6_, s_81__5_, s_81__4_, 
        s_81__3_, s_81__2_, s_81__1_, s_81__0_}) );
  reg_7 R8 ( .Reset(n1298), .Clk(Clk), .Load(n2), .Din({s_67__31_, s_67__30_, 
        s_67__29_, s_67__28_, s_67__27_, s_67__26_, s_67__25_, s_67__24_, 
        s_67__23_, s_67__22_, s_67__21_, s_67__20_, s_67__19_, s_67__18_, 
        s_67__17_, s_67__16_, s_67__15_, s_67__14_, s_67__13_, s_67__12_, 
        s_67__11_, s_67__10_, s_67__9_, s_67__8_, s_67__7_, s_67__6_, s_67__5_, 
        s_67__4_, s_67__3_, s_67__2_, s_67__1_, s_67__0_}), .Dout(sr[223:192])
         );
  reg_6 R9 ( .Reset(n1293), .Clk(Clk), .Load(n2), .Din({s_66__31_, s_66__30_, 
        s_66__29_, s_66__28_, s_66__27_, s_66__26_, s_66__25_, s_66__24_, 
        s_66__23_, s_66__22_, s_66__21_, s_66__20_, s_66__19_, s_66__18_, 
        s_66__17_, s_66__16_, s_66__15_, s_66__14_, s_66__13_, s_66__12_, 
        s_66__11_, s_66__10_, s_66__9_, s_66__8_, s_66__7_, s_66__6_, s_66__5_, 
        s_66__4_, s_66__3_, s_66__2_, s_66__1_, s_66__0_}), .Dout(sr[191:160])
         );
  adder_23 S80 ( .A(sr[223:192]), .B(sr[191:160]), .O({s_80__31_, s_80__30_, 
        s_80__29_, s_80__28_, s_80__27_, s_80__26_, s_80__25_, s_80__24_, 
        s_80__23_, s_80__22_, s_80__21_, s_80__20_, s_80__19_, s_80__18_, 
        s_80__17_, s_80__16_, s_80__15_, s_80__14_, s_80__13_, s_80__12_, 
        s_80__11_, s_80__10_, s_80__9_, s_80__8_, s_80__7_, s_80__6_, s_80__5_, 
        s_80__4_, s_80__3_, s_80__2_, s_80__1_, s_80__0_}) );
  adder_22 S67 ( .A({s_63__31_, s_63__30_, s_63__29_, s_63__28_, s_63__27_, 
        s_63__26_, s_63__25_, s_63__24_, s_63__23_, s_63__22_, s_63__21_, 
        s_63__20_, s_63__19_, s_63__18_, s_63__17_, s_63__16_, s_63__15_, 
        s_63__14_, s_63__13_, s_63__12_, s_63__11_, s_63__10_, s_63__9_, 
        s_63__8_, s_63__7_, s_63__6_, s_63__5_, s_63__4_, s_63__3_, s_63__2_, 
        s_63__1_, s_63__0_}), .B({s_62__31_, s_62__30_, s_62__29_, s_62__28_, 
        s_62__27_, s_62__26_, s_62__25_, s_62__24_, s_62__23_, s_62__22_, 
        s_62__21_, s_62__20_, s_62__19_, s_62__18_, s_62__17_, s_62__16_, 
        s_62__15_, s_62__14_, s_62__13_, s_62__12_, s_62__11_, s_62__10_, 
        s_62__9_, s_62__8_, s_62__7_, s_62__6_, s_62__5_, s_62__4_, s_62__3_, 
        s_62__2_, s_62__1_, s_62__0_}), .O({s_67__31_, s_67__30_, s_67__29_, 
        s_67__28_, s_67__27_, s_67__26_, s_67__25_, s_67__24_, s_67__23_, 
        s_67__22_, s_67__21_, s_67__20_, s_67__19_, s_67__18_, s_67__17_, 
        s_67__16_, s_67__15_, s_67__14_, s_67__13_, s_67__12_, s_67__11_, 
        s_67__10_, s_67__9_, s_67__8_, s_67__7_, s_67__6_, s_67__5_, s_67__4_, 
        s_67__3_, s_67__2_, s_67__1_, s_67__0_}) );
  adder_21 S63 ( .A({y_2__29_, y_2__28_, y_2__27_, y_2__26_, y_2__25_, 
        y_2__24_, y_2__23_, y_2__22_, n1291, n1289, n1285, n1283, n1281, n1278, 
        n1276, n1273, n1270, n1267, n1264, n1260, n1257, n1255, n1253, n1250, 
        n1247, n1244, n1241, n1238, n1234, n1232, n1, n1}), .B({y_2__22_, 
        n1291, n1288, n1285, n1283, n1281, n1279, n1275, n1272, n1269, n1267, 
        n1264, n1261, n1258, n1255, n1252, n1249, n1246, n1243, n1241, n1237, 
        n1234, n1232, n1, n1, n1, n1, n1, n1, n1, n1, n1}), .O({s_63__31_, 
        s_63__30_, s_63__29_, s_63__28_, s_63__27_, s_63__26_, s_63__25_, 
        s_63__24_, s_63__23_, s_63__22_, s_63__21_, s_63__20_, s_63__19_, 
        s_63__18_, s_63__17_, s_63__16_, s_63__15_, s_63__14_, s_63__13_, 
        s_63__12_, s_63__11_, s_63__10_, s_63__9_, s_63__8_, s_63__7_, 
        s_63__6_, s_63__5_, s_63__4_, s_63__3_, s_63__2_, s_63__1_, s_63__0_})
         );
  adder_20 S62 ( .A({Input[284:256], n1, n1, n1}), .B({Input[283:256], n1, n1, 
        n1, n1}), .O({s_62__31_, s_62__30_, s_62__29_, s_62__28_, s_62__27_, 
        s_62__26_, s_62__25_, s_62__24_, s_62__23_, s_62__22_, s_62__21_, 
        s_62__20_, s_62__19_, s_62__18_, s_62__17_, s_62__16_, s_62__15_, 
        s_62__14_, s_62__13_, s_62__12_, s_62__11_, s_62__10_, s_62__9_, 
        s_62__8_, s_62__7_, s_62__6_, s_62__5_, s_62__4_, s_62__3_, s_62__2_, 
        s_62__1_, s_62__0_}) );
  adder_19 S66 ( .A({s_65__31_, s_65__30_, s_65__29_, s_65__28_, s_65__27_, 
        s_65__26_, s_65__25_, s_65__24_, s_65__23_, s_65__22_, s_65__21_, 
        s_65__20_, s_65__19_, s_65__18_, s_65__17_, s_65__16_, s_65__15_, 
        s_65__14_, s_65__13_, s_65__12_, s_65__11_, s_65__10_, s_65__9_, 
        s_65__8_, s_65__7_, s_65__6_, s_65__5_, s_65__4_, s_65__3_, s_65__2_, 
        s_65__1_, s_65__0_}), .B({s_64__31_, s_64__30_, s_64__29_, s_64__28_, 
        s_64__27_, s_64__26_, s_64__25_, s_64__24_, s_64__23_, s_64__22_, 
        s_64__21_, s_64__20_, s_64__19_, s_64__18_, s_64__17_, s_64__16_, 
        s_64__15_, s_64__14_, s_64__13_, s_64__12_, s_64__11_, s_64__10_, 
        s_64__9_, s_64__8_, s_64__7_, s_64__6_, s_64__5_, s_64__4_, s_64__3_, 
        s_64__2_, s_64__1_, s_64__0_}), .O({s_66__31_, s_66__30_, s_66__29_, 
        s_66__28_, s_66__27_, s_66__26_, s_66__25_, s_66__24_, s_66__23_, 
        s_66__22_, s_66__21_, s_66__20_, s_66__19_, s_66__18_, s_66__17_, 
        s_66__16_, s_66__15_, s_66__14_, s_66__13_, s_66__12_, s_66__11_, 
        s_66__10_, s_66__9_, s_66__8_, s_66__7_, s_66__6_, s_66__5_, s_66__4_, 
        s_66__3_, s_66__2_, s_66__1_, s_66__0_}) );
  adder_18 S65 ( .A({Input[318:288], n1}), .B({y_1__31_, y_1__30_, y_1__29_, 
        y_1__28_, y_1__27_, y_1__26_, y_1__25_, y_1__24_, y_1__23_, y_1__22_, 
        n1181, y_1__20_, n1184, n1183, n1198, n1215, n1203, n1214, n1211, 
        n1209, n1222, y_1__10_, n1225, n1218, n1229, n1188, n1228, n1217, 
        n1226, n1220, n1213, n1189}), .O({s_65__31_, s_65__30_, s_65__29_, 
        s_65__28_, s_65__27_, s_65__26_, s_65__25_, s_65__24_, s_65__23_, 
        s_65__22_, s_65__21_, s_65__20_, s_65__19_, s_65__18_, s_65__17_, 
        s_65__16_, s_65__15_, s_65__14_, s_65__13_, s_65__12_, s_65__11_, 
        s_65__10_, s_65__9_, s_65__8_, s_65__7_, s_65__6_, s_65__5_, s_65__4_, 
        s_65__3_, s_65__2_, s_65__1_, s_65__0_}) );
  adder_17 S64 ( .A({n1292, n1289, n1286, n1283, n1281, n1279, n1275, n1273, 
        n1270, n1266, n1263, n1261, n1258, n1255, n1252, n1250, n1247, n1244, 
        n1240, n1238, n1235, n1232, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1}), 
        .B(Input[319:288]), .O({s_64__31_, s_64__30_, s_64__29_, s_64__28_, 
        s_64__27_, s_64__26_, s_64__25_, s_64__24_, s_64__23_, s_64__22_, 
        s_64__21_, s_64__20_, s_64__19_, s_64__18_, s_64__17_, s_64__16_, 
        s_64__15_, s_64__14_, s_64__13_, s_64__12_, s_64__11_, s_64__10_, 
        s_64__9_, s_64__8_, s_64__7_, s_64__6_, s_64__5_, s_64__4_, s_64__3_, 
        s_64__2_, s_64__1_, s_64__0_}) );
  reg_5 R10 ( .Reset(n1293), .Clk(Clk), .Load(n2), .Din({s_69__31_, s_69__30_, 
        s_69__29_, s_69__28_, s_69__27_, s_69__26_, s_69__25_, s_69__24_, 
        s_69__23_, s_69__22_, s_69__21_, s_69__20_, s_69__19_, s_69__18_, 
        s_69__17_, s_69__16_, s_69__15_, s_69__14_, s_69__13_, s_69__12_, 
        s_69__11_, s_69__10_, s_69__9_, s_69__8_, s_69__7_, s_69__6_, s_69__5_, 
        s_69__4_, s_69__3_, s_69__2_, s_69__1_, s_69__0_}), .Dout(sr[159:128])
         );
  reg_4 R11 ( .Reset(n1295), .Clk(Clk), .Load(n2), .Din({s_68__31_, s_68__30_, 
        s_68__29_, s_68__28_, s_68__27_, s_68__26_, s_68__25_, s_68__24_, 
        s_68__23_, s_68__22_, s_68__21_, s_68__20_, s_68__19_, s_68__18_, 
        s_68__17_, s_68__16_, s_68__15_, s_68__14_, s_68__13_, s_68__12_, 
        s_68__11_, s_68__10_, s_68__9_, s_68__8_, s_68__7_, s_68__6_, s_68__5_, 
        s_68__4_, s_68__3_, s_68__2_, s_68__1_, s_68__0_}), .Dout(sr[127:96])
         );
  adder_16 S79 ( .A(sr[159:128]), .B(sr[127:96]), .O({s_79__31_, s_79__30_, 
        s_79__29_, s_79__28_, s_79__27_, s_79__26_, s_79__25_, s_79__24_, 
        s_79__23_, s_79__22_, s_79__21_, s_79__20_, s_79__19_, s_79__18_, 
        s_79__17_, s_79__16_, s_79__15_, s_79__14_, s_79__13_, s_79__12_, 
        s_79__11_, s_79__10_, s_79__9_, s_79__8_, s_79__7_, s_79__6_, s_79__5_, 
        s_79__4_, s_79__3_, s_79__2_, s_79__1_, s_79__0_}) );
  adder_15 S69 ( .A({s_59__31_, s_59__30_, s_59__29_, s_59__28_, s_59__27_, 
        s_59__26_, s_59__25_, s_59__24_, s_59__23_, s_59__22_, s_59__21_, 
        s_59__20_, s_59__19_, s_59__18_, s_59__17_, s_59__16_, s_59__15_, 
        s_59__14_, s_59__13_, s_59__12_, s_59__11_, s_59__10_, s_59__9_, 
        s_59__8_, s_59__7_, s_59__6_, s_59__5_, s_59__4_, s_59__3_, s_59__2_, 
        s_59__1_, s_59__0_}), .B({s_58__31_, s_58__30_, s_58__29_, s_58__28_, 
        s_58__27_, s_58__26_, s_58__25_, s_58__24_, s_58__23_, s_58__22_, 
        s_58__21_, s_58__20_, s_58__19_, s_58__18_, s_58__17_, s_58__16_, 
        s_58__15_, s_58__14_, s_58__13_, s_58__12_, s_58__11_, s_58__10_, 
        s_58__9_, s_58__8_, s_58__7_, s_58__6_, s_58__5_, s_58__4_, s_58__3_, 
        s_58__2_, s_58__1_, s_58__0_}), .O({s_69__31_, s_69__30_, s_69__29_, 
        s_69__28_, s_69__27_, s_69__26_, s_69__25_, s_69__24_, s_69__23_, 
        s_69__22_, s_69__21_, s_69__20_, s_69__19_, s_69__18_, s_69__17_, 
        s_69__16_, s_69__15_, s_69__14_, s_69__13_, s_69__12_, s_69__11_, 
        s_69__10_, s_69__9_, s_69__8_, s_69__7_, s_69__6_, s_69__5_, s_69__4_, 
        s_69__3_, s_69__2_, s_69__1_, s_69__0_}) );
  adder_14 S59 ( .A({Input[250:224], n1, n1, n1, n1, n1}), .B({Input[249:224], 
        n1, n1, n1, n1, n1, n1}), .O({s_59__31_, s_59__30_, s_59__29_, 
        s_59__28_, s_59__27_, s_59__26_, s_59__25_, s_59__24_, s_59__23_, 
        s_59__22_, s_59__21_, s_59__20_, s_59__19_, s_59__18_, s_59__17_, 
        s_59__16_, s_59__15_, s_59__14_, s_59__13_, s_59__12_, s_59__11_, 
        s_59__10_, s_59__9_, s_59__8_, s_59__7_, s_59__6_, s_59__5_, s_59__4_, 
        s_59__3_, s_59__2_, s_59__1_, s_59__0_}) );
  adder_13 S58 ( .A({y_4__28_, y_4__27_, y_4__26_, y_4__25_, y_4__24_, 
        y_4__23_, y_4__22_, y_4__21_, y_4__20_, y_4__19_, y_4__18_, y_4__17_, 
        y_4__16_, y_4__15_, y_4__14_, n1201, y_4__12_, n1196, y_4__10_, 
        y_4__9_, n1180, y_4__7_, y_4__6_, y_4__5_, n1182, y_4__3_, y_4__2_, 
        y_4__1_, y_4__0_, n1, n1, n1}), .B({y_4__25_, y_4__24_, y_4__23_, 
        y_4__22_, y_4__21_, y_4__20_, y_4__19_, y_4__18_, y_4__17_, y_4__16_, 
        y_4__15_, y_4__14_, y_4__13_, y_4__12_, n1196, y_4__10_, y_4__9_, 
        n1180, y_4__7_, y_4__6_, y_4__5_, n1182, y_4__3_, y_4__2_, y_4__1_, 
        y_4__0_, n1, n1, n1, n1, n1, n1}), .O({s_58__31_, s_58__30_, s_58__29_, 
        s_58__28_, s_58__27_, s_58__26_, s_58__25_, s_58__24_, s_58__23_, 
        s_58__22_, s_58__21_, s_58__20_, s_58__19_, s_58__18_, s_58__17_, 
        s_58__16_, s_58__15_, s_58__14_, s_58__13_, s_58__12_, s_58__11_, 
        s_58__10_, s_58__9_, s_58__8_, s_58__7_, s_58__6_, s_58__5_, s_58__4_, 
        s_58__3_, s_58__2_, s_58__1_, s_58__0_}) );
  adder_12 S68 ( .A({s_61__31_, s_61__30_, s_61__29_, s_61__28_, s_61__27_, 
        s_61__26_, s_61__25_, s_61__24_, s_61__23_, s_61__22_, s_61__21_, 
        s_61__20_, s_61__19_, s_61__18_, s_61__17_, s_61__16_, s_61__15_, 
        s_61__14_, s_61__13_, s_61__12_, s_61__11_, s_61__10_, s_61__9_, 
        s_61__8_, s_61__7_, s_61__6_, s_61__5_, s_61__4_, s_61__3_, s_61__2_, 
        s_61__1_, s_61__0_}), .B({s_60__31_, s_60__30_, s_60__29_, s_60__28_, 
        s_60__27_, s_60__26_, s_60__25_, s_60__24_, s_60__23_, s_60__22_, 
        s_60__21_, s_60__20_, s_60__19_, s_60__18_, s_60__17_, s_60__16_, 
        s_60__15_, s_60__14_, s_60__13_, s_60__12_, s_60__11_, s_60__10_, 
        s_60__9_, s_60__8_, s_60__7_, s_60__6_, s_60__5_, s_60__4_, s_60__3_, 
        s_60__2_, s_60__1_, s_60__0_}), .O({s_68__31_, s_68__30_, s_68__29_, 
        s_68__28_, s_68__27_, s_68__26_, s_68__25_, s_68__24_, s_68__23_, 
        s_68__22_, s_68__21_, s_68__20_, s_68__19_, s_68__18_, s_68__17_, 
        s_68__16_, s_68__15_, s_68__14_, s_68__13_, s_68__12_, s_68__11_, 
        s_68__10_, s_68__9_, s_68__8_, s_68__7_, s_68__6_, s_68__5_, s_68__4_, 
        s_68__3_, s_68__2_, s_68__1_, s_68__0_}) );
  adder_11 S61 ( .A({y_3__23_, y_3__22_, y_3__21_, y_3__20_, y_3__19_, 
        y_3__18_, y_3__17_, y_3__16_, y_3__15_, y_3__14_, n1200, y_3__12_, 
        n1187, y_3__10_, y_3__9_, y_3__8_, y_3__7_, y_3__6_, y_3__5_, y_3__4_, 
        y_3__3_, y_3__2_, y_3__1_, y_3__0_, n1, n1, n1, n1, n1, n1, n1, n1}), 
        .B(Input[287:256]), .O({s_61__31_, s_61__30_, s_61__29_, s_61__28_, 
        s_61__27_, s_61__26_, s_61__25_, s_61__24_, s_61__23_, s_61__22_, 
        s_61__21_, s_61__20_, s_61__19_, s_61__18_, s_61__17_, s_61__16_, 
        s_61__15_, s_61__14_, s_61__13_, s_61__12_, s_61__11_, s_61__10_, 
        s_61__9_, s_61__8_, s_61__7_, s_61__6_, s_61__5_, s_61__4_, s_61__3_, 
        s_61__2_, s_61__1_, s_61__0_}) );
  adder_10 S60 ( .A({y_3__31_, y_3__30_, y_3__29_, y_3__28_, y_3__27_, 
        y_3__26_, y_3__25_, y_3__24_, y_3__23_, y_3__22_, y_3__21_, y_3__20_, 
        y_3__19_, y_3__18_, y_3__17_, y_3__16_, y_3__15_, y_3__14_, n1200, 
        y_3__12_, n1187, y_3__10_, y_3__9_, y_3__8_, y_3__7_, y_3__6_, y_3__5_, 
        y_3__4_, y_3__3_, y_3__2_, y_3__1_, y_3__0_}), .B({y_3__25_, y_3__24_, 
        y_3__23_, y_3__22_, y_3__21_, y_3__20_, y_3__19_, y_3__18_, y_3__17_, 
        y_3__16_, y_3__15_, y_3__14_, n1200, y_3__12_, n1187, y_3__10_, 
        y_3__9_, y_3__8_, y_3__7_, y_3__6_, y_3__5_, y_3__4_, y_3__3_, y_3__2_, 
        y_3__1_, y_3__0_, n1, n1, n1, n1, n1, n1}), .O({s_60__31_, s_60__30_, 
        s_60__29_, s_60__28_, s_60__27_, s_60__26_, s_60__25_, s_60__24_, 
        s_60__23_, s_60__22_, s_60__21_, s_60__20_, s_60__19_, s_60__18_, 
        s_60__17_, s_60__16_, s_60__15_, s_60__14_, s_60__13_, s_60__12_, 
        s_60__11_, s_60__10_, s_60__9_, s_60__8_, s_60__7_, s_60__6_, s_60__5_, 
        s_60__4_, s_60__3_, s_60__2_, s_60__1_, s_60__0_}) );
  reg_3 R12 ( .Reset(n1297), .Clk(Clk), .Load(n2), .Din({s_83__31_, s_83__30_, 
        s_83__29_, s_83__28_, s_83__27_, s_83__26_, s_83__25_, s_83__24_, 
        s_83__23_, s_83__22_, s_83__21_, s_83__20_, s_83__19_, s_83__18_, 
        s_83__17_, s_83__16_, s_83__15_, s_83__14_, s_83__13_, s_83__12_, 
        s_83__11_, s_83__10_, s_83__9_, s_83__8_, s_83__7_, s_83__6_, s_83__5_, 
        s_83__4_, s_83__3_, s_83__2_, s_83__1_, s_83__0_}), .Dout(sr[95:64])
         );
  adder_9 S86 ( .A({y_1__26_, y_1__25_, y_1__24_, y_1__23_, y_1__22_, n1181, 
        y_1__20_, n1184, n1183, n1198, n1215, n1203, n1214, n1211, n1209, 
        n1222, y_1__10_, n1225, n1218, y_1__7_, n1224, n1228, n1217, n1226, 
        n1220, n1213, y_1__0_, n1, n1, n1, n1, n1}), .B(sr[95:64]), .O({
        s_86__31_, s_86__30_, s_86__29_, s_86__28_, s_86__27_, s_86__26_, 
        s_86__25_, s_86__24_, s_86__23_, s_86__22_, s_86__21_, s_86__20_, 
        s_86__19_, s_86__18_, s_86__17_, s_86__16_, s_86__15_, s_86__14_, 
        s_86__13_, s_86__12_, s_86__11_, s_86__10_, s_86__9_, s_86__8_, 
        s_86__7_, s_86__6_, s_86__5_, s_86__4_, s_86__3_, s_86__2_, s_86__1_, 
        s_86__0_}) );
  adder_8 S83 ( .A({s_76__31_, s_76__30_, s_76__29_, s_76__28_, s_76__27_, 
        s_76__26_, s_76__25_, s_76__24_, s_76__23_, s_76__22_, s_76__21_, 
        s_76__20_, s_76__19_, s_76__18_, s_76__17_, s_76__16_, s_76__15_, 
        s_76__14_, s_76__13_, s_76__12_, s_76__11_, s_76__10_, s_76__9_, 
        s_76__8_, s_76__7_, s_76__6_, s_76__5_, s_76__4_, s_76__3_, s_76__2_, 
        s_76__1_, s_76__0_}), .B({s_75__31_, s_75__30_, s_75__29_, s_75__28_, 
        s_75__27_, s_75__26_, s_75__25_, s_75__24_, s_75__23_, s_75__22_, 
        s_75__21_, s_75__20_, s_75__19_, s_75__18_, s_75__17_, s_75__16_, 
        s_75__15_, s_75__14_, s_75__13_, s_75__12_, s_75__11_, s_75__10_, 
        s_75__9_, s_75__8_, s_75__7_, s_75__6_, s_75__5_, s_75__4_, s_75__3_, 
        s_75__2_, s_75__1_, s_75__0_}), .O({s_83__31_, s_83__30_, s_83__29_, 
        s_83__28_, s_83__27_, s_83__26_, s_83__25_, s_83__24_, s_83__23_, 
        s_83__22_, s_83__21_, s_83__20_, s_83__19_, s_83__18_, s_83__17_, 
        s_83__16_, s_83__15_, s_83__14_, s_83__13_, s_83__12_, s_83__11_, 
        s_83__10_, s_83__9_, s_83__8_, s_83__7_, s_83__6_, s_83__5_, s_83__4_, 
        s_83__3_, s_83__2_, s_83__1_, s_83__0_}) );
  reg_2 R13 ( .Reset(n1293), .Clk(Clk), .Load(n2), .Din({s_47__31_, s_47__30_, 
        s_47__29_, s_47__28_, s_47__27_, s_47__26_, s_47__25_, s_47__24_, 
        s_47__23_, s_47__22_, s_47__21_, s_47__20_, s_47__19_, s_47__18_, 
        s_47__17_, s_47__16_, s_47__15_, s_47__14_, s_47__13_, s_47__12_, 
        s_47__11_, s_47__10_, s_47__9_, s_47__8_, s_47__7_, s_47__6_, s_47__5_, 
        s_47__4_, s_47__3_, s_47__2_, s_47__1_, s_47__0_}), .Dout(sr[63:32])
         );
  reg_1 R14 ( .Reset(n1294), .Clk(Clk), .Load(n2), .Din({s_74__31_, s_74__30_, 
        s_74__29_, s_74__28_, s_74__27_, s_74__26_, s_74__25_, s_74__24_, 
        s_74__23_, s_74__22_, s_74__21_, s_74__20_, s_74__19_, s_74__18_, 
        s_74__17_, s_74__16_, s_74__15_, s_74__14_, s_74__13_, s_74__12_, 
        s_74__11_, s_74__10_, s_74__9_, s_74__8_, s_74__7_, s_74__6_, s_74__5_, 
        s_74__4_, s_74__3_, s_74__2_, s_74__1_, s_74__0_}), .Dout(sr[31:0]) );
  adder_7 S76 ( .A(sr[63:32]), .B(sr[31:0]), .O({s_76__31_, s_76__30_, 
        s_76__29_, s_76__28_, s_76__27_, s_76__26_, s_76__25_, s_76__24_, 
        s_76__23_, s_76__22_, s_76__21_, s_76__20_, s_76__19_, s_76__18_, 
        s_76__17_, s_76__16_, s_76__15_, s_76__14_, s_76__13_, s_76__12_, 
        s_76__11_, s_76__10_, s_76__9_, s_76__8_, s_76__7_, s_76__6_, s_76__5_, 
        s_76__4_, s_76__3_, s_76__2_, s_76__1_, s_76__0_}) );
  adder_6 S47 ( .A(Input[31:0]), .B({Input[30:0], n1}), .O({s_47__31_, 
        s_47__30_, s_47__29_, s_47__28_, s_47__27_, s_47__26_, s_47__25_, 
        s_47__24_, s_47__23_, s_47__22_, s_47__21_, s_47__20_, s_47__19_, 
        s_47__18_, s_47__17_, s_47__16_, s_47__15_, s_47__14_, s_47__13_, 
        s_47__12_, s_47__11_, s_47__10_, s_47__9_, s_47__8_, s_47__7_, 
        s_47__6_, s_47__5_, s_47__4_, s_47__3_, s_47__2_, s_47__1_, s_47__0_})
         );
  adder_5 S74 ( .A({s_49__31_, s_49__30_, s_49__29_, s_49__28_, s_49__27_, 
        s_49__26_, s_49__25_, s_49__24_, s_49__23_, s_49__22_, s_49__21_, 
        s_49__20_, s_49__19_, s_49__18_, s_49__17_, s_49__16_, s_49__15_, 
        s_49__14_, s_49__13_, s_49__12_, s_49__11_, s_49__10_, s_49__9_, 
        s_49__8_, s_49__7_, s_49__6_, s_49__5_, s_49__4_, s_49__3_, s_49__2_, 
        s_49__1_, s_49__0_}), .B({s_48__31_, s_48__30_, s_48__29_, s_48__28_, 
        s_48__27_, s_48__26_, s_48__25_, s_48__24_, s_48__23_, s_48__22_, 
        s_48__21_, s_48__20_, s_48__19_, s_48__18_, s_48__17_, s_48__16_, 
        s_48__15_, s_48__14_, s_48__13_, s_48__12_, s_48__11_, s_48__10_, 
        s_48__9_, s_48__8_, s_48__7_, s_48__6_, s_48__5_, s_48__4_, s_48__3_, 
        s_48__2_, s_48__1_, s_48__0_}), .O({s_74__31_, s_74__30_, s_74__29_, 
        s_74__28_, s_74__27_, s_74__26_, s_74__25_, s_74__24_, s_74__23_, 
        s_74__22_, s_74__21_, s_74__20_, s_74__19_, s_74__18_, s_74__17_, 
        s_74__16_, s_74__15_, s_74__14_, s_74__13_, s_74__12_, s_74__11_, 
        s_74__10_, s_74__9_, s_74__8_, s_74__7_, s_74__6_, s_74__5_, s_74__4_, 
        s_74__3_, s_74__2_, s_74__1_, s_74__0_}) );
  adder_4 S49 ( .A({Input[59:39], n1207, n1191, n1205, Input[35:32], n1, n1, 
        n1, n1}), .B({Input[90:68], n1193, Input[66:64], n1, n1, n1, n1, n1}), 
        .O({s_49__31_, s_49__30_, s_49__29_, s_49__28_, s_49__27_, s_49__26_, 
        s_49__25_, s_49__24_, s_49__23_, s_49__22_, s_49__21_, s_49__20_, 
        s_49__19_, s_49__18_, s_49__17_, s_49__16_, s_49__15_, s_49__14_, 
        s_49__13_, s_49__12_, s_49__11_, s_49__10_, s_49__9_, s_49__8_, 
        s_49__7_, s_49__6_, s_49__5_, s_49__4_, s_49__3_, s_49__2_, s_49__1_, 
        s_49__0_}) );
  adder_3 S48 ( .A({Input[63:39], n1207, n1191, n1205, Input[35], n1208, n1185, 
        Input[32]}), .B({Input[60:39], n1207, n1191, n1205, Input[35:32], n1, 
        n1, n1}), .O({s_48__31_, s_48__30_, s_48__29_, s_48__28_, s_48__27_, 
        s_48__26_, s_48__25_, s_48__24_, s_48__23_, s_48__22_, s_48__21_, 
        s_48__20_, s_48__19_, s_48__18_, s_48__17_, s_48__16_, s_48__15_, 
        s_48__14_, s_48__13_, s_48__12_, s_48__11_, s_48__10_, s_48__9_, 
        s_48__8_, s_48__7_, s_48__6_, s_48__5_, s_48__4_, s_48__3_, s_48__2_, 
        s_48__1_, s_48__0_}) );
  adder_2 S75 ( .A({y_2__25_, y_2__24_, y_2__23_, y_2__22_, n1292, n1288, 
        n1285, n1283, n1281, n1278, n1276, n1272, n1269, n1266, n1264, n1261, 
        n1257, n1255, n1253, n1249, n1246, n1243, n1241, n1237, n1234, n1232, 
        n1, n1, n1, n1, n1, n1}), .B({y_2__23_, y_2__22_, n1291, n1288, n1286, 
        n1283, n1281, n1279, n1275, n1273, n1269, n1266, n1263, n1260, n1258, 
        n1255, n1252, n1249, n1246, n1243, n1240, n1237, n1235, n1232, n1, n1, 
        n1, n1, n1, n1, n1, n1}), .O({s_75__31_, s_75__30_, s_75__29_, 
        s_75__28_, s_75__27_, s_75__26_, s_75__25_, s_75__24_, s_75__23_, 
        s_75__22_, s_75__21_, s_75__20_, s_75__19_, s_75__18_, s_75__17_, 
        s_75__16_, s_75__15_, s_75__14_, s_75__13_, s_75__12_, s_75__11_, 
        s_75__10_, s_75__9_, s_75__8_, s_75__7_, s_75__6_, s_75__5_, s_75__4_, 
        s_75__3_, s_75__2_, s_75__1_, s_75__0_}) );
  adder_1 S90 ( .A({y_1__31_, y_1__30_, y_1__29_, y_1__28_, y_1__27_, y_1__26_, 
        y_1__25_, y_1__24_, y_1__23_, y_1__22_, n1181, y_1__20_, n1184, n1183, 
        n1198, n1215, n1203, n1214, n1211, n1209, n1222, y_1__10_, n1225, 
        n1218, n1229, n1188, n1228, n1217, n1226, n1220, n1213, n1189}), .B({
        y_1__29_, y_1__28_, y_1__27_, y_1__26_, y_1__25_, y_1__24_, y_1__23_, 
        y_1__22_, n1181, y_1__20_, n1184, n1183, n1198, n1215, n1203, n1214, 
        n1211, n1209, n1222, y_1__10_, n1225, n1218, n1229, n1224, n1228, 
        n1217, n1226, n1220, n1213, y_1__0_, n1, n1}), .O({s_90__31_, 
        s_90__30_, s_90__29_, s_90__28_, s_90__27_, s_90__26_, s_90__25_, 
        s_90__24_, s_90__23_, s_90__22_, s_90__21_, s_90__20_, s_90__19_, 
        s_90__18_, s_90__17_, s_90__16_, s_90__15_, s_90__14_, s_90__13_, 
        s_90__12_, s_90__11_, s_90__10_, s_90__9_, s_90__8_, s_90__7_, 
        s_90__6_, s_90__5_, s_90__4_, s_90__3_, s_90__2_, s_90__1_, s_90__0_})
         );
  BUF8 U3 ( .A(y_4__13_), .Q(n1201) );
  INV12 U4 ( .A(n1265), .Q(n1266) );
  CLKIN8 U5 ( .A(y_2__12_), .Q(n1265) );
  CLKIN15 U6 ( .A(n1204), .Q(n1205) );
  INV12 U7 ( .A(n1262), .Q(n1264) );
  INV6 U8 ( .A(y_5__9_), .Q(n1177) );
  INV10 U9 ( .A(n1177), .Q(n1178) );
  INV4 U10 ( .A(n1277), .Q(n1279) );
  INV8 U11 ( .A(n1268), .Q(n1269) );
  CLKIN12 U12 ( .A(n1274), .Q(n1276) );
  INV15 U13 ( .A(n1242), .Q(n1243) );
  INV8 U14 ( .A(n1268), .Q(n1270) );
  INV15 U15 ( .A(n1248), .Q(n1249) );
  INV15 U16 ( .A(n1202), .Q(n1203) );
  CLKIN6 U17 ( .A(Input[38]), .Q(n1206) );
  CLKIN15 U18 ( .A(n1230), .Q(n1232) );
  INV12 U19 ( .A(n1197), .Q(n1198) );
  CLKIN12 U20 ( .A(y_2__15_), .Q(n1274) );
  INV6 U21 ( .A(y_1__1_), .Q(n1212) );
  BUF15 U22 ( .A(y_1__7_), .Q(n1229) );
  INV15 U23 ( .A(n1216), .Q(n1217) );
  CLKIN15 U24 ( .A(n1239), .Q(n1240) );
  INV15 U25 ( .A(n1239), .Q(n1241) );
  INV10 U26 ( .A(y_2__3_), .Q(n1239) );
  INV15 U27 ( .A(n1190), .Q(n1191) );
  CLKIN12 U28 ( .A(y_2__10_), .Q(n1259) );
  INV12 U29 ( .A(n1259), .Q(n1261) );
  INV12 U30 ( .A(y_2__5_), .Q(n1245) );
  INV6 U31 ( .A(y_2__16_), .Q(n1277) );
  INV15 U32 ( .A(n1248), .Q(n1250) );
  CLKIN12 U33 ( .A(y_2__6_), .Q(n1248) );
  INV15 U34 ( .A(n1256), .Q(n1258) );
  CLKIN12 U35 ( .A(n1274), .Q(n1275) );
  INV15 U36 ( .A(n1210), .Q(n1211) );
  INV8 U37 ( .A(y_4__8_), .Q(n1179) );
  INV15 U38 ( .A(n1179), .Q(n1180) );
  CLKIN6 U39 ( .A(n1277), .Q(n1278) );
  INV15 U40 ( .A(n1245), .Q(n1246) );
  CLKIN12 U41 ( .A(y_2__4_), .Q(n1242) );
  INV15 U42 ( .A(n1236), .Q(n1237) );
  INV15 U43 ( .A(n1282), .Q(n1283) );
  CLKIN15 U44 ( .A(n1262), .Q(n1263) );
  INV10 U45 ( .A(y_2__11_), .Q(n1262) );
  INV10 U46 ( .A(y_2__13_), .Q(n1268) );
  CLKIN6 U47 ( .A(n1284), .Q(n1286) );
  CLKIN6 U48 ( .A(y_2__19_), .Q(n1284) );
  INV12 U49 ( .A(n1230), .Q(n1231) );
  CLKIN12 U50 ( .A(y_2__0_), .Q(n1230) );
  CLKBU15 U51 ( .A(y_1__9_), .Q(n1225) );
  CLKBU15 U52 ( .A(y_1__14_), .Q(n1214) );
  INV15 U53 ( .A(n1233), .Q(n1235) );
  INV12 U54 ( .A(n1265), .Q(n1267) );
  INV12 U55 ( .A(n1256), .Q(n1257) );
  INV12 U56 ( .A(n1192), .Q(n1193) );
  INV6 U57 ( .A(n1287), .Q(n1288) );
  CLKIN8 U58 ( .A(y_2__9_), .Q(n1256) );
  CLKIN6 U59 ( .A(y_2__14_), .Q(n1271) );
  CLKIN8 U60 ( .A(y_2__1_), .Q(n1233) );
  INV8 U61 ( .A(y_2__2_), .Q(n1236) );
  CLKIN6 U62 ( .A(y_2__18_), .Q(n1282) );
  INV3 U63 ( .A(y_2__21_), .Q(n1290) );
  INV8 U64 ( .A(y_1__6_), .Q(n1223) );
  INV12 U65 ( .A(n1245), .Q(n1247) );
  INV8 U66 ( .A(n1284), .Q(n1285) );
  INV6 U67 ( .A(n1287), .Q(n1289) );
  INV3 U68 ( .A(y_1__17_), .Q(n1197) );
  INV12 U69 ( .A(n1271), .Q(n1272) );
  INV6 U70 ( .A(n1290), .Q(n1291) );
  INV10 U71 ( .A(n1223), .Q(n1188) );
  INV12 U72 ( .A(n1223), .Q(n1224) );
  BUF8 U73 ( .A(y_1__21_), .Q(n1181) );
  BUF15 U74 ( .A(y_4__4_), .Q(n1182) );
  INV6 U75 ( .A(y_2__17_), .Q(n1280) );
  INV12 U76 ( .A(n1280), .Q(n1281) );
  BUF6 U77 ( .A(y_1__18_), .Q(n1183) );
  BUF8 U78 ( .A(y_1__19_), .Q(n1184) );
  CLKIN12 U79 ( .A(n1242), .Q(n1244) );
  INV6 U80 ( .A(y_1__5_), .Q(n1227) );
  BUF2 U81 ( .A(Input[33]), .Q(n1185) );
  BUF15 U82 ( .A(y_1__16_), .Q(n1215) );
  CLKIN12 U83 ( .A(n1233), .Q(n1234) );
  CLKIN6 U84 ( .A(y_3__11_), .Q(n1186) );
  INV12 U85 ( .A(n1186), .Q(n1187) );
  INV15 U86 ( .A(n1219), .Q(n1220) );
  INV6 U87 ( .A(y_1__2_), .Q(n1219) );
  CLKBU2 U88 ( .A(y_1__0_), .Q(n1189) );
  INV6 U89 ( .A(Input[37]), .Q(n1190) );
  CLKIN15 U90 ( .A(n1212), .Q(n1213) );
  BUF15 U91 ( .A(y_1__8_), .Q(n1218) );
  BUF15 U92 ( .A(y_1__12_), .Q(n1209) );
  INV12 U93 ( .A(n1206), .Q(n1207) );
  BUF15 U94 ( .A(y_1__3_), .Q(n1226) );
  INV6 U95 ( .A(Input[67]), .Q(n1192) );
  INV6 U96 ( .A(Input[36]), .Q(n1204) );
  INV6 U97 ( .A(y_2__8_), .Q(n1254) );
  INV15 U98 ( .A(n1254), .Q(n1255) );
  INV15 U99 ( .A(n1221), .Q(n1222) );
  BUF2 U100 ( .A(y_4__5_), .Q(n1194) );
  INV12 U101 ( .A(n1236), .Q(n1238) );
  CLKIN6 U102 ( .A(y_4__11_), .Q(n1195) );
  INV12 U103 ( .A(n1195), .Q(n1196) );
  CLKIN6 U104 ( .A(y_3__13_), .Q(n1199) );
  INV12 U105 ( .A(n1199), .Q(n1200) );
  INV15 U106 ( .A(n1227), .Q(n1228) );
  CLKIN12 U107 ( .A(y_2__7_), .Q(n1251) );
  CLKIN6 U108 ( .A(y_1__15_), .Q(n1202) );
  INV15 U109 ( .A(n1251), .Q(n1252) );
  BUF2 U110 ( .A(Input[34]), .Q(n1208) );
  INV15 U111 ( .A(n1251), .Q(n1253) );
  INV15 U112 ( .A(n1259), .Q(n1260) );
  INV12 U113 ( .A(n1271), .Q(n1273) );
  INV6 U114 ( .A(n1290), .Q(n1292) );
  INV3 U115 ( .A(n1296), .Q(n1299) );
  INV3 U116 ( .A(n1296), .Q(n1298) );
  INV3 U117 ( .A(n1296), .Q(n1297) );
  CLKBU2 U118 ( .A(n1300), .Q(n1295) );
  CLKBU2 U119 ( .A(n1300), .Q(n1294) );
  CLKBU2 U120 ( .A(n1300), .Q(n1293) );
  CLKIN6 U121 ( .A(y_2__20_), .Q(n1287) );
  CLKIN6 U122 ( .A(y_1__4_), .Q(n1216) );
  INV3 U123 ( .A(n1300), .Q(n1296) );
  CLKBU2 U124 ( .A(Reset), .Q(n1300) );
  LOGIC1 U125 ( .Q(n2) );
  LOGIC0 U126 ( .Q(n1) );
  CLKIN6 U127 ( .A(y_1__13_), .Q(n1210) );
  CLKIN6 U128 ( .A(y_1__11_), .Q(n1221) );
endmodule


module reg_25 ( Reset, Clk, Load, Din, Dout );
  input [31:0] Din;
  output [31:0] Dout;
  input Reset, Clk, Load;
  wire   n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32,
         n35, n47, n49, n51, n53, n55, n57, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n125, n126,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407;

  DF3 Dout_reg_1_ ( .D(n112), .C(Clk), .Q(Dout[1]), .QN(n100) );
  DF3 Dout_reg_0_ ( .D(n113), .C(Clk), .Q(Dout[0]), .QN(n102) );
  DF3 Dout_reg_2_ ( .D(n111), .C(Clk), .Q(Dout[2]), .QN(n101) );
  DF3 Dout_reg_3_ ( .D(n110), .C(Clk), .Q(Dout[3]), .QN(n95) );
  DF3 Dout_reg_6_ ( .D(n107), .C(Clk), .Q(Dout[6]), .QN(n98) );
  DF3 Dout_reg_5_ ( .D(n108), .C(Clk), .Q(Dout[5]), .QN(n97) );
  DF3 Dout_reg_8_ ( .D(n105), .C(Clk), .Q(Dout[8]), .QN(n93) );
  OAI222 U3 ( .A(n6), .B(n372), .C(n374), .D(n396), .Q(n83) );
  OAI222 U4 ( .A(n8), .B(n372), .C(n373), .D(n395), .Q(n82) );
  OAI222 U5 ( .A(n10), .B(n372), .C(n125), .D(n394), .Q(n81) );
  OAI222 U6 ( .A(n12), .B(n372), .C(n374), .D(n393), .Q(n80) );
  OAI222 U7 ( .A(n14), .B(n372), .C(n373), .D(n392), .Q(n79) );
  OAI222 U8 ( .A(n16), .B(n372), .C(n125), .D(n378), .Q(n78) );
  OAI222 U9 ( .A(n18), .B(n372), .C(n374), .D(n391), .Q(n77) );
  OAI222 U10 ( .A(n20), .B(n372), .C(n373), .D(n376), .Q(n76) );
  OAI222 U11 ( .A(n22), .B(n372), .C(n125), .D(n377), .Q(n75) );
  OAI222 U12 ( .A(n24), .B(n372), .C(n382), .D(n374), .Q(n74) );
  OAI222 U13 ( .A(n26), .B(n372), .C(n373), .D(n381), .Q(n73) );
  OAI222 U14 ( .A(n28), .B(n372), .C(n125), .D(n379), .Q(n72) );
  OAI222 U15 ( .A(n30), .B(n372), .C(n374), .D(n380), .Q(n71) );
  OAI222 U16 ( .A(n32), .B(n372), .C(n373), .D(n383), .Q(n70) );
  OAI222 U17 ( .A(n35), .B(n372), .C(n385), .D(n125), .Q(n69) );
  OAI222 U18 ( .A(n47), .B(n372), .C(n387), .D(n374), .Q(n68) );
  OAI222 U19 ( .A(n49), .B(n372), .C(n373), .D(n384), .Q(n67) );
  OAI222 U20 ( .A(n51), .B(n372), .C(n125), .D(n386), .Q(n66) );
  OAI222 U21 ( .A(n53), .B(n372), .C(n390), .D(n374), .Q(n65) );
  OAI222 U22 ( .A(n55), .B(n372), .C(n373), .D(n389), .Q(n64) );
  OAI222 U23 ( .A(n57), .B(n372), .C(n125), .D(n388), .Q(n63) );
  OAI222 U24 ( .A(n102), .B(n372), .C(n374), .D(n407), .Q(n113) );
  OAI222 U25 ( .A(n100), .B(n372), .C(n373), .D(n406), .Q(n112) );
  OAI222 U26 ( .A(n101), .B(n372), .C(n125), .D(n405), .Q(n111) );
  OAI222 U27 ( .A(n95), .B(n372), .C(n374), .D(n404), .Q(n110) );
  OAI222 U28 ( .A(n96), .B(n372), .C(n373), .D(n403), .Q(n109) );
  OAI222 U29 ( .A(n97), .B(n372), .C(n125), .D(n402), .Q(n108) );
  OAI222 U30 ( .A(n98), .B(n372), .C(n374), .D(n401), .Q(n107) );
  OAI222 U31 ( .A(n99), .B(n372), .C(n373), .D(n400), .Q(n106) );
  OAI222 U32 ( .A(n93), .B(n372), .C(n125), .D(n398), .Q(n105) );
  OAI222 U33 ( .A(n92), .B(n372), .C(n374), .D(n399), .Q(n104) );
  OAI222 U34 ( .A(n94), .B(n372), .C(n373), .D(n397), .Q(n103) );
  DF1 Dout_reg_20_ ( .D(n74), .C(Clk), .Q(Dout[20]), .QN(n24) );
  DF1 Dout_reg_29_ ( .D(n65), .C(Clk), .Q(Dout[29]), .QN(n53) );
  DF1 Dout_reg_22_ ( .D(n72), .C(Clk), .Q(Dout[22]), .QN(n28) );
  DF1 Dout_reg_19_ ( .D(n75), .C(Clk), .Q(Dout[19]), .QN(n22) );
  DF1 Dout_reg_23_ ( .D(n71), .C(Clk), .Q(Dout[23]), .QN(n30) );
  DF1 Dout_reg_26_ ( .D(n68), .C(Clk), .Q(Dout[26]), .QN(n47) );
  DF1 Dout_reg_31_ ( .D(n63), .C(Clk), .Q(Dout[31]), .QN(n57) );
  DF1 Dout_reg_17_ ( .D(n77), .C(Clk), .Q(Dout[17]), .QN(n18) );
  DF1 Dout_reg_28_ ( .D(n66), .C(Clk), .Q(Dout[28]), .QN(n51) );
  DF1 Dout_reg_27_ ( .D(n67), .C(Clk), .Q(Dout[27]), .QN(n49) );
  DF1 Dout_reg_25_ ( .D(n69), .C(Clk), .Q(Dout[25]), .QN(n35) );
  DF1 Dout_reg_24_ ( .D(n70), .C(Clk), .Q(Dout[24]), .QN(n32) );
  DF1 Dout_reg_4_ ( .D(n109), .C(Clk), .Q(Dout[4]), .QN(n96) );
  DF1 Dout_reg_16_ ( .D(n78), .C(Clk), .Q(Dout[16]), .QN(n16) );
  DF1 Dout_reg_10_ ( .D(n103), .C(Clk), .Q(Dout[10]), .QN(n94) );
  DF1 Dout_reg_9_ ( .D(n104), .C(Clk), .Q(Dout[9]), .QN(n92) );
  DF1 Dout_reg_15_ ( .D(n79), .C(Clk), .Q(Dout[15]), .QN(n14) );
  DF1 Dout_reg_21_ ( .D(n73), .C(Clk), .Q(Dout[21]), .QN(n26) );
  DF1 Dout_reg_13_ ( .D(n81), .C(Clk), .Q(Dout[13]), .QN(n10) );
  DF1 Dout_reg_11_ ( .D(n83), .C(Clk), .Q(Dout[11]), .QN(n6) );
  DF1 Dout_reg_14_ ( .D(n80), .C(Clk), .Q(Dout[14]), .QN(n12) );
  DF1 Dout_reg_12_ ( .D(n82), .C(Clk), .Q(Dout[12]), .QN(n8) );
  DF1 Dout_reg_7_ ( .D(n106), .C(Clk), .Q(Dout[7]), .QN(n99) );
  DF1 Dout_reg_18_ ( .D(n76), .C(Clk), .Q(Dout[18]), .QN(n20) );
  DF1 Dout_reg_30_ ( .D(n64), .C(Clk), .Q(Dout[30]), .QN(n55) );
  INV3 U35 ( .A(Din[17]), .Q(n391) );
  INV2 U36 ( .A(Din[20]), .Q(n382) );
  INV3 U37 ( .A(Din[30]), .Q(n389) );
  INV3 U38 ( .A(Din[31]), .Q(n388) );
  CLKIN3 U39 ( .A(Din[6]), .Q(n401) );
  INV2 U40 ( .A(Din[4]), .Q(n403) );
  INV2 U41 ( .A(Din[16]), .Q(n378) );
  INV2 U42 ( .A(Din[8]), .Q(n398) );
  CLKIN3 U43 ( .A(Din[5]), .Q(n402) );
  NAND22 U44 ( .A(n375), .B(n372), .Q(n374) );
  NAND22 U45 ( .A(n375), .B(n372), .Q(n373) );
  NAND22 U46 ( .A(n375), .B(n372), .Q(n125) );
  INV3 U47 ( .A(n126), .Q(n372) );
  INV3 U48 ( .A(Din[29]), .Q(n390) );
  INV3 U49 ( .A(Din[23]), .Q(n380) );
  INV3 U50 ( .A(Din[9]), .Q(n399) );
  INV3 U51 ( .A(Din[12]), .Q(n395) );
  INV3 U52 ( .A(Din[14]), .Q(n393) );
  INV3 U53 ( .A(Din[11]), .Q(n396) );
  INV3 U54 ( .A(Din[15]), .Q(n392) );
  INV3 U55 ( .A(Din[10]), .Q(n397) );
  INV3 U56 ( .A(Din[7]), .Q(n400) );
  INV3 U57 ( .A(Din[1]), .Q(n406) );
  INV3 U58 ( .A(Din[19]), .Q(n377) );
  INV3 U59 ( .A(Din[22]), .Q(n379) );
  INV3 U60 ( .A(Din[13]), .Q(n394) );
  INV3 U61 ( .A(Din[2]), .Q(n405) );
  INV3 U62 ( .A(Din[3]), .Q(n404) );
  INV3 U63 ( .A(Din[0]), .Q(n407) );
  NOR20 U64 ( .A(Load), .B(Reset), .Q(n126) );
  INV3 U65 ( .A(Reset), .Q(n375) );
  INV3 U66 ( .A(Din[21]), .Q(n381) );
  INV3 U67 ( .A(Din[18]), .Q(n376) );
  INV3 U68 ( .A(Din[24]), .Q(n383) );
  INV3 U69 ( .A(Din[26]), .Q(n387) );
  INV3 U70 ( .A(Din[28]), .Q(n386) );
  INV3 U71 ( .A(Din[25]), .Q(n385) );
  INV3 U72 ( .A(Din[27]), .Q(n384) );
endmodule


module iir_sol_wrapper ( Reset, Clk, Input, Output );
  input [31:0] Input;
  output [31:0] Output;
  input Reset, Clk;
  wire   del_1__31_, del_1__30_, del_1__29_, del_1__28_, del_1__27_,
         del_1__26_, del_1__25_, del_1__24_, del_1__23_, del_1__22_,
         del_1__21_, del_1__20_, del_1__19_, del_1__18_, del_1__17_,
         del_1__16_, del_1__15_, del_1__14_, del_1__13_, del_1__12_,
         del_1__11_, del_1__10_, del_1__9_, del_1__8_, del_1__7_, del_1__6_,
         del_1__5_, del_1__4_, del_1__3_, del_1__2_, del_1__1_, del_1__0_,
         del_2__31_, del_2__30_, del_2__29_, del_2__28_, del_2__27_,
         del_2__26_, del_2__25_, del_2__24_, del_2__23_, del_2__22_,
         del_2__21_, del_2__20_, del_2__19_, del_2__18_, del_2__17_,
         del_2__16_, del_2__15_, del_2__14_, del_2__13_, del_2__12_,
         del_2__11_, del_2__10_, del_2__9_, del_2__8_, del_2__7_, del_2__6_,
         del_2__5_, del_2__4_, del_2__3_, del_2__2_, del_2__1_, del_2__0_,
         del_3__31_, del_3__30_, del_3__29_, del_3__28_, del_3__27_,
         del_3__26_, del_3__25_, del_3__24_, del_3__23_, del_3__22_,
         del_3__21_, del_3__20_, del_3__19_, del_3__18_, del_3__17_,
         del_3__16_, del_3__15_, del_3__14_, del_3__13_, del_3__12_,
         del_3__11_, del_3__10_, del_3__9_, del_3__8_, del_3__7_, del_3__6_,
         del_3__5_, del_3__4_, del_3__3_, del_3__2_, del_3__1_, del_3__0_,
         del_4__31_, del_4__30_, del_4__29_, del_4__28_, del_4__27_,
         del_4__26_, del_4__25_, del_4__24_, del_4__23_, del_4__22_,
         del_4__21_, del_4__20_, del_4__19_, del_4__18_, del_4__17_,
         del_4__16_, del_4__15_, del_4__14_, del_4__13_, del_4__12_,
         del_4__11_, del_4__10_, del_4__9_, del_4__8_, del_4__7_, del_4__6_,
         del_4__5_, del_4__4_, del_4__3_, del_4__2_, del_4__1_, del_4__0_,
         del_5__31_, del_5__30_, del_5__29_, del_5__28_, del_5__27_,
         del_5__26_, del_5__25_, del_5__24_, del_5__23_, del_5__22_,
         del_5__21_, del_5__20_, del_5__19_, del_5__18_, del_5__17_,
         del_5__16_, del_5__15_, del_5__14_, del_5__13_, del_5__12_,
         del_5__11_, del_5__10_, del_5__9_, del_5__8_, del_5__7_, del_5__6_,
         del_5__5_, del_5__4_, del_5__3_, del_5__2_, del_5__1_, del_5__0_,
         del_6__31_, del_6__30_, del_6__29_, del_6__28_, del_6__27_,
         del_6__26_, del_6__25_, del_6__24_, del_6__23_, del_6__22_,
         del_6__21_, del_6__20_, del_6__19_, del_6__18_, del_6__17_,
         del_6__16_, del_6__15_, del_6__14_, del_6__13_, del_6__12_,
         del_6__11_, del_6__10_, del_6__9_, del_6__8_, del_6__7_, del_6__6_,
         del_6__5_, del_6__4_, del_6__3_, del_6__2_, del_6__1_, del_6__0_,
         del_7__31_, del_7__30_, del_7__29_, del_7__28_, del_7__27_,
         del_7__26_, del_7__25_, del_7__24_, del_7__23_, del_7__22_,
         del_7__21_, del_7__20_, del_7__19_, del_7__18_, del_7__17_,
         del_7__16_, del_7__15_, del_7__14_, del_7__13_, del_7__12_,
         del_7__11_, del_7__10_, del_7__9_, del_7__8_, del_7__7_, del_7__6_,
         del_7__5_, del_7__4_, del_7__3_, del_7__2_, del_7__1_, del_7__0_,
         del_8__31_, del_8__30_, del_8__29_, del_8__28_, del_8__27_,
         del_8__26_, del_8__25_, del_8__24_, del_8__23_, del_8__22_,
         del_8__21_, del_8__20_, del_8__19_, del_8__18_, del_8__17_,
         del_8__16_, del_8__15_, del_8__14_, del_8__13_, del_8__12_,
         del_8__11_, del_8__10_, del_8__9_, del_8__8_, del_8__7_, del_8__6_,
         del_8__5_, del_8__4_, del_8__3_, del_8__2_, del_8__1_, del_8__0_,
         del_9__31_, del_9__30_, del_9__29_, del_9__28_, del_9__27_,
         del_9__26_, del_9__25_, del_9__24_, del_9__23_, del_9__22_,
         del_9__21_, del_9__20_, del_9__19_, del_9__18_, del_9__17_,
         del_9__16_, del_9__15_, del_9__14_, del_9__13_, del_9__12_,
         del_9__11_, del_9__10_, del_9__9_, del_9__8_, del_9__7_, del_9__6_,
         del_9__5_, del_9__4_, del_9__3_, del_9__2_, del_9__1_, del_9__0_,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283;
  wire   [31:0] outs;

  reg_0 R_0 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din(Input), .Dout({
        del_1__31_, del_1__30_, del_1__29_, del_1__28_, del_1__27_, del_1__26_, 
        del_1__25_, del_1__24_, del_1__23_, del_1__22_, del_1__21_, del_1__20_, 
        del_1__19_, del_1__18_, del_1__17_, del_1__16_, del_1__15_, del_1__14_, 
        del_1__13_, del_1__12_, del_1__11_, del_1__10_, del_1__9_, del_1__8_, 
        del_1__7_, del_1__6_, del_1__5_, del_1__4_, del_1__3_, del_1__2_, 
        del_1__1_, del_1__0_}) );
  reg_33 R_1 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din({del_1__31_, 
        del_1__30_, del_1__29_, del_1__28_, del_1__27_, del_1__26_, del_1__25_, 
        del_1__24_, del_1__23_, del_1__22_, del_1__21_, del_1__20_, del_1__19_, 
        del_1__18_, del_1__17_, del_1__16_, del_1__15_, del_1__14_, del_1__13_, 
        del_1__12_, del_1__11_, n274, n281, del_1__8_, del_1__7_, del_1__6_, 
        n273, del_1__4_, del_1__3_, del_1__2_, del_1__1_, del_1__0_}), .Dout({
        del_2__31_, del_2__30_, del_2__29_, del_2__28_, del_2__27_, del_2__26_, 
        del_2__25_, del_2__24_, del_2__23_, del_2__22_, del_2__21_, del_2__20_, 
        del_2__19_, del_2__18_, del_2__17_, del_2__16_, del_2__15_, del_2__14_, 
        del_2__13_, del_2__12_, del_2__11_, del_2__10_, del_2__9_, del_2__8_, 
        del_2__7_, del_2__6_, del_2__5_, del_2__4_, del_2__3_, del_2__2_, 
        del_2__1_, del_2__0_}) );
  reg_32 R_2 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din({del_2__31_, 
        del_2__30_, del_2__29_, del_2__28_, del_2__27_, del_2__26_, del_2__25_, 
        del_2__24_, del_2__23_, del_2__22_, del_2__21_, del_2__20_, del_2__19_, 
        del_2__18_, del_2__17_, del_2__16_, del_2__15_, del_2__14_, del_2__13_, 
        del_2__12_, del_2__11_, del_2__10_, del_2__9_, del_2__8_, del_2__7_, 
        del_2__6_, del_2__5_, del_2__4_, del_2__3_, del_2__2_, del_2__1_, 
        del_2__0_}), .Dout({del_3__31_, del_3__30_, del_3__29_, del_3__28_, 
        del_3__27_, del_3__26_, del_3__25_, del_3__24_, del_3__23_, del_3__22_, 
        del_3__21_, del_3__20_, del_3__19_, del_3__18_, del_3__17_, del_3__16_, 
        del_3__15_, del_3__14_, del_3__13_, del_3__12_, del_3__11_, del_3__10_, 
        del_3__9_, del_3__8_, del_3__7_, del_3__6_, del_3__5_, del_3__4_, 
        del_3__3_, del_3__2_, del_3__1_, del_3__0_}) );
  reg_31 R_3 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din({del_3__31_, 
        del_3__30_, del_3__29_, del_3__28_, del_3__27_, del_3__26_, del_3__25_, 
        del_3__24_, del_3__23_, del_3__22_, del_3__21_, del_3__20_, del_3__19_, 
        del_3__18_, del_3__17_, del_3__16_, del_3__15_, del_3__14_, del_3__13_, 
        del_3__12_, del_3__11_, del_3__10_, del_3__9_, del_3__8_, del_3__7_, 
        del_3__6_, del_3__5_, del_3__4_, del_3__3_, del_3__2_, del_3__1_, 
        del_3__0_}), .Dout({del_4__31_, del_4__30_, del_4__29_, del_4__28_, 
        del_4__27_, del_4__26_, del_4__25_, del_4__24_, del_4__23_, del_4__22_, 
        del_4__21_, del_4__20_, del_4__19_, del_4__18_, del_4__17_, del_4__16_, 
        del_4__15_, del_4__14_, del_4__13_, del_4__12_, del_4__11_, del_4__10_, 
        del_4__9_, del_4__8_, del_4__7_, del_4__6_, del_4__5_, del_4__4_, 
        del_4__3_, del_4__2_, del_4__1_, del_4__0_}) );
  reg_30 R_4 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din({del_4__31_, 
        del_4__30_, del_4__29_, del_4__28_, del_4__27_, del_4__26_, del_4__25_, 
        del_4__24_, del_4__23_, del_4__22_, del_4__21_, del_4__20_, del_4__19_, 
        del_4__18_, del_4__17_, del_4__16_, del_4__15_, del_4__14_, del_4__13_, 
        del_4__12_, del_4__11_, del_4__10_, del_4__9_, del_4__8_, del_4__7_, 
        n277, del_4__5_, del_4__4_, del_4__3_, del_4__2_, del_4__1_, del_4__0_}), .Dout({del_5__31_, del_5__30_, del_5__29_, del_5__28_, del_5__27_, 
        del_5__26_, del_5__25_, del_5__24_, del_5__23_, del_5__22_, del_5__21_, 
        del_5__20_, del_5__19_, del_5__18_, del_5__17_, del_5__16_, del_5__15_, 
        del_5__14_, del_5__13_, del_5__12_, del_5__11_, del_5__10_, del_5__9_, 
        del_5__8_, del_5__7_, del_5__6_, del_5__5_, del_5__4_, del_5__3_, 
        del_5__2_, del_5__1_, del_5__0_}) );
  reg_29 R_5 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din({del_5__31_, 
        del_5__30_, del_5__29_, del_5__28_, del_5__27_, del_5__26_, del_5__25_, 
        del_5__24_, del_5__23_, del_5__22_, del_5__21_, del_5__20_, del_5__19_, 
        del_5__18_, del_5__17_, del_5__16_, del_5__15_, del_5__14_, del_5__13_, 
        del_5__12_, del_5__11_, del_5__10_, del_5__9_, del_5__8_, del_5__7_, 
        del_5__6_, del_5__5_, del_5__4_, del_5__3_, del_5__2_, del_5__1_, 
        del_5__0_}), .Dout({del_6__31_, del_6__30_, del_6__29_, del_6__28_, 
        del_6__27_, del_6__26_, del_6__25_, del_6__24_, del_6__23_, del_6__22_, 
        del_6__21_, del_6__20_, del_6__19_, del_6__18_, del_6__17_, del_6__16_, 
        del_6__15_, del_6__14_, del_6__13_, del_6__12_, del_6__11_, del_6__10_, 
        del_6__9_, del_6__8_, del_6__7_, del_6__6_, del_6__5_, del_6__4_, 
        del_6__3_, del_6__2_, del_6__1_, del_6__0_}) );
  reg_28 R_6 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din({del_6__31_, 
        del_6__30_, del_6__29_, del_6__28_, del_6__27_, del_6__26_, del_6__25_, 
        del_6__24_, del_6__23_, del_6__22_, del_6__21_, del_6__20_, del_6__19_, 
        del_6__18_, del_6__17_, del_6__16_, del_6__15_, del_6__14_, del_6__13_, 
        del_6__12_, del_6__11_, del_6__10_, del_6__9_, del_6__8_, del_6__7_, 
        del_6__6_, del_6__5_, del_6__4_, del_6__3_, del_6__2_, del_6__1_, 
        del_6__0_}), .Dout({del_7__31_, del_7__30_, del_7__29_, del_7__28_, 
        del_7__27_, del_7__26_, del_7__25_, del_7__24_, del_7__23_, del_7__22_, 
        del_7__21_, del_7__20_, del_7__19_, del_7__18_, del_7__17_, del_7__16_, 
        del_7__15_, del_7__14_, del_7__13_, del_7__12_, del_7__11_, del_7__10_, 
        del_7__9_, del_7__8_, del_7__7_, del_7__6_, del_7__5_, del_7__4_, 
        del_7__3_, del_7__2_, del_7__1_, del_7__0_}) );
  reg_27 R_7 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din({del_7__31_, 
        del_7__30_, del_7__29_, del_7__28_, del_7__27_, del_7__26_, del_7__25_, 
        del_7__24_, del_7__23_, del_7__22_, del_7__21_, del_7__20_, del_7__19_, 
        del_7__18_, del_7__17_, del_7__16_, del_7__15_, del_7__14_, del_7__13_, 
        del_7__12_, del_7__11_, del_7__10_, del_7__9_, del_7__8_, del_7__7_, 
        del_7__6_, del_7__5_, del_7__4_, del_7__3_, del_7__2_, del_7__1_, 
        del_7__0_}), .Dout({del_8__31_, del_8__30_, del_8__29_, del_8__28_, 
        del_8__27_, del_8__26_, del_8__25_, del_8__24_, del_8__23_, del_8__22_, 
        del_8__21_, del_8__20_, del_8__19_, del_8__18_, del_8__17_, del_8__16_, 
        del_8__15_, del_8__14_, del_8__13_, del_8__12_, del_8__11_, del_8__10_, 
        del_8__9_, del_8__8_, del_8__7_, del_8__6_, del_8__5_, del_8__4_, 
        del_8__3_, del_8__2_, del_8__1_, del_8__0_}) );
  reg_26 R_8 ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din({del_8__31_, 
        del_8__30_, del_8__29_, del_8__28_, del_8__27_, del_8__26_, del_8__25_, 
        del_8__24_, del_8__23_, del_8__22_, del_8__21_, del_8__20_, del_8__19_, 
        del_8__18_, del_8__17_, del_8__16_, del_8__15_, del_8__14_, del_8__13_, 
        del_8__12_, del_8__11_, n279, del_8__9_, n283, del_8__7_, del_8__6_, 
        del_8__5_, n275, del_8__3_, del_8__2_, del_8__1_, del_8__0_}), .Dout({
        del_9__31_, del_9__30_, del_9__29_, del_9__28_, del_9__27_, del_9__26_, 
        del_9__25_, del_9__24_, del_9__23_, del_9__22_, del_9__21_, del_9__20_, 
        del_9__19_, del_9__18_, del_9__17_, del_9__16_, del_9__15_, del_9__14_, 
        del_9__13_, del_9__12_, del_9__11_, del_9__10_, del_9__9_, del_9__8_, 
        del_9__7_, del_9__6_, del_9__5_, del_9__4_, del_9__3_, del_9__2_, 
        del_9__1_, del_9__0_}) );
  iir_sol U1 ( .Reset(Reset), .Clk(Clk), .Input({Input, del_1__31_, del_1__30_, 
        del_1__29_, del_1__28_, del_1__27_, del_1__26_, del_1__25_, del_1__24_, 
        del_1__23_, del_1__22_, del_1__21_, del_1__20_, del_1__19_, del_1__18_, 
        del_1__17_, del_1__16_, del_1__15_, del_1__14_, del_1__13_, del_1__12_, 
        del_1__11_, del_1__10_, n281, del_1__8_, del_1__7_, del_1__6_, 
        del_1__5_, del_1__4_, del_1__3_, del_1__2_, del_1__1_, del_1__0_, 
        del_2__31_, del_2__30_, del_2__29_, del_2__28_, del_2__27_, del_2__26_, 
        del_2__25_, del_2__24_, del_2__23_, del_2__22_, del_2__21_, del_2__20_, 
        del_2__19_, del_2__18_, del_2__17_, del_2__16_, del_2__15_, del_2__14_, 
        del_2__13_, del_2__12_, del_2__11_, del_2__10_, del_2__9_, del_2__8_, 
        del_2__7_, del_2__6_, del_2__5_, del_2__4_, del_2__3_, del_2__2_, 
        del_2__1_, del_2__0_, del_3__31_, del_3__30_, del_3__29_, del_3__28_, 
        del_3__27_, del_3__26_, del_3__25_, del_3__24_, del_3__23_, del_3__22_, 
        del_3__21_, del_3__20_, del_3__19_, del_3__18_, del_3__17_, del_3__16_, 
        del_3__15_, del_3__14_, del_3__13_, del_3__12_, del_3__11_, del_3__10_, 
        del_3__9_, del_3__8_, del_3__7_, del_3__6_, del_3__5_, del_3__4_, 
        del_3__3_, del_3__2_, del_3__1_, del_3__0_, del_4__31_, del_4__30_, 
        del_4__29_, del_4__28_, del_4__27_, del_4__26_, del_4__25_, del_4__24_, 
        del_4__23_, del_4__22_, del_4__21_, del_4__20_, del_4__19_, del_4__18_, 
        del_4__17_, del_4__16_, del_4__15_, del_4__14_, del_4__13_, del_4__12_, 
        del_4__11_, del_4__10_, del_4__9_, del_4__8_, del_4__7_, n277, 
        del_4__5_, del_4__4_, del_4__3_, del_4__2_, del_4__1_, del_4__0_, 
        del_5__31_, del_5__30_, del_5__29_, del_5__28_, del_5__27_, del_5__26_, 
        del_5__25_, del_5__24_, del_5__23_, del_5__22_, del_5__21_, del_5__20_, 
        del_5__19_, del_5__18_, del_5__17_, del_5__16_, del_5__15_, del_5__14_, 
        del_5__13_, del_5__12_, del_5__11_, del_5__10_, del_5__9_, del_5__8_, 
        del_5__7_, del_5__6_, del_5__5_, del_5__4_, del_5__3_, del_5__2_, 
        del_5__1_, del_5__0_, del_6__31_, del_6__30_, del_6__29_, del_6__28_, 
        del_6__27_, del_6__26_, del_6__25_, del_6__24_, del_6__23_, del_6__22_, 
        del_6__21_, del_6__20_, del_6__19_, del_6__18_, del_6__17_, del_6__16_, 
        del_6__15_, del_6__14_, del_6__13_, del_6__12_, del_6__11_, del_6__10_, 
        del_6__9_, del_6__8_, del_6__7_, del_6__6_, del_6__5_, del_6__4_, 
        del_6__3_, del_6__2_, del_6__1_, del_6__0_, del_7__31_, del_7__30_, 
        del_7__29_, del_7__28_, del_7__27_, del_7__26_, del_7__25_, del_7__24_, 
        del_7__23_, del_7__22_, del_7__21_, del_7__20_, del_7__19_, del_7__18_, 
        del_7__17_, del_7__16_, del_7__15_, del_7__14_, del_7__13_, del_7__12_, 
        del_7__11_, del_7__10_, del_7__9_, del_7__8_, del_7__7_, del_7__6_, 
        del_7__5_, del_7__4_, del_7__3_, del_7__2_, del_7__1_, del_7__0_, 
        del_8__31_, del_8__30_, del_8__29_, del_8__28_, del_8__27_, del_8__26_, 
        del_8__25_, del_8__24_, del_8__23_, del_8__22_, del_8__21_, del_8__20_, 
        del_8__19_, del_8__18_, del_8__17_, del_8__16_, del_8__15_, del_8__14_, 
        del_8__13_, del_8__12_, del_8__11_, n279, del_8__9_, n283, del_8__7_, 
        del_8__6_, del_8__5_, del_8__4_, del_8__3_, del_8__2_, del_8__1_, 
        del_8__0_, del_9__31_, del_9__30_, del_9__29_, del_9__28_, del_9__27_, 
        del_9__26_, del_9__25_, del_9__24_, del_9__23_, del_9__22_, del_9__21_, 
        del_9__20_, del_9__19_, del_9__18_, del_9__17_, del_9__16_, del_9__15_, 
        del_9__14_, del_9__13_, del_9__12_, del_9__11_, del_9__10_, del_9__9_, 
        del_9__8_, del_9__7_, del_9__6_, del_9__5_, del_9__4_, del_9__3_, 
        del_9__2_, del_9__1_, del_9__0_}), .Output(outs) );
  reg_25 R_o ( .Reset(Reset), .Clk(Clk), .Load(n272), .Din(outs), .Dout(Output) );
  INV12 U11 ( .A(n276), .Q(n277) );
  BUF2 U12 ( .A(del_1__5_), .Q(n273) );
  INV15 U13 ( .A(n280), .Q(n281) );
  BUF2 U14 ( .A(del_1__10_), .Q(n274) );
  BUF2 U15 ( .A(del_8__4_), .Q(n275) );
  CLKIN6 U16 ( .A(del_4__6_), .Q(n276) );
  CLKIN6 U17 ( .A(del_8__10_), .Q(n278) );
  INV12 U18 ( .A(n278), .Q(n279) );
  CLKIN6 U19 ( .A(del_1__9_), .Q(n280) );
  INV6 U20 ( .A(del_8__8_), .Q(n282) );
  INV12 U21 ( .A(n282), .Q(n283) );
  LOGIC1 U22 ( .Q(n272) );
endmodule

